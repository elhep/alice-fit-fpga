----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:22:33 08/05/2016 
-- Design Name: 
-- Module Name:    fit - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
library UNISIM;
use UNISIM.vcomponents.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.all;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

library work;
use work.PM12_pkg.all;

use work.fit_gbt_common_package.all;
use work.fit_gbt_board_package.all;

entity PM12 is
  port
  (
    TDCCLK1_P : in std_logic;
    TDCCLK1_N : in std_logic;
    RDA1_P    : in std_logic;
    RDA1_N    : in std_logic;
    RSA1_P    : in std_logic;
    RSA1_N    : in std_logic;
    RDB1_P    : in std_logic;
    RDB1_N    : in std_logic;
    RSB1_P    : in std_logic;
    RSB1_N    : in std_logic;
    RDC1_P    : in std_logic;
    RDC1_N    : in std_logic;
    RSC1_P    : in std_logic;
    RSC1_N    : in std_logic;
    RDD1_P    : in std_logic;
    RDD1_N    : in std_logic;
    RSD1_P    : in std_logic;
    RSD1_N    : in std_logic;
    INA1_P    : in std_logic;
    INA1_N    : in std_logic;
    INB1_P    : in std_logic;
    INB1_N    : in std_logic;
    INC1_P    : in std_logic;
    INC1_N    : in std_logic;
    IND1_P    : in std_logic;
    IND1_N    : in std_logic;
    DI1       : in std_logic_vector (12 downto 0);
    DI2       : in std_logic_vector (12 downto 0);
    DI3       : in std_logic_vector (12 downto 0);
    DI4       : in std_logic_vector (12 downto 0);
    STR1      : in std_logic;
    STR2      : in std_logic;
    STR3      : in std_logic;
    STR4      : in std_logic;
    MCLK1_P   : in std_logic;
    MCLK1_N   : in std_logic;

    TDCCLK2_P : in std_logic;
    TDCCLK2_N : in std_logic;
    RDA2_P    : in std_logic;
    RDA2_N    : in std_logic;
    RSA2_P    : in std_logic;
    RSA2_N    : in std_logic;
    RDB2_P    : in std_logic;
    RDB2_N    : in std_logic;
    RSB2_P    : in std_logic;
    RSB2_N    : in std_logic;
    RDC2_P    : in std_logic;
    RDC2_N    : in std_logic;
    RSC2_P    : in std_logic;
    RSC2_N    : in std_logic;
    RDD2_P    : in std_logic;
    RDD2_N    : in std_logic;
    RSD2_P    : in std_logic;
    RSD2_N    : in std_logic;
    INA2_P    : in std_logic;
    INA2_N    : in std_logic;
    INB2_P    : in std_logic;
    INB2_N    : in std_logic;
    INC2_P    : in std_logic;
    INC2_N    : in std_logic;
    IND2_P    : in std_logic;
    IND2_N    : in std_logic;
    DI5       : in std_logic_vector (12 downto 0);
    DI6       : in std_logic_vector (12 downto 0);
    DI7       : in std_logic_vector (12 downto 0);
    DI8       : in std_logic_vector (12 downto 0);
    STR5      : in std_logic;
    STR6      : in std_logic;
    STR7      : in std_logic;
    STR8      : in std_logic;
    MCLK2_P   : in std_logic;
    MCLK2_N   : in std_logic;

    TDCCLK3_P : in std_logic;
    TDCCLK3_N : in std_logic;
    RDA3_P    : in std_logic;
    RDA3_N    : in std_logic;
    RSA3_P    : in std_logic;
    RSA3_N    : in std_logic;
    RDB3_P    : in std_logic;
    RDB3_N    : in std_logic;
    RSB3_P    : in std_logic;
    RSB3_N    : in std_logic;
    RDC3_P    : in std_logic;
    RDC3_N    : in std_logic;
    RSC3_P    : in std_logic;
    RSC3_N    : in std_logic;
    RDD3_P    : in std_logic;
    RDD3_N    : in std_logic;
    RSD3_P    : in std_logic;
    RSD3_N    : in std_logic;
    INA3_P    : in std_logic;
    INA3_N    : in std_logic;
    INB3_P    : in std_logic;
    INB3_N    : in std_logic;
    INC3_P    : in std_logic;
    INC3_N    : in std_logic;
    IND3_P    : in std_logic;
    IND3_N    : in std_logic;
    DI9       : in std_logic_vector (12 downto 0);
    DI10      : in std_logic_vector (12 downto 0);
    DI11      : in std_logic_vector (12 downto 0);
    DI12      : in std_logic_vector (12 downto 0);
    STR9      : in std_logic;
    STR10     : in std_logic;
    STR11     : in std_logic;
    STR12     : in std_logic;
    MCLK3_P   : in std_logic;
    MCLK3_N   : in std_logic;

    SCK       : in std_logic;
    MISO      : out std_logic;
    MOSI      : in std_logic;
    CS        : in std_logic;

    RST       : in std_logic;
    IRQ       : out std_logic;

    AT0_P     : out std_logic;
    AT0_N     : out std_logic;
    AT1_P     : out std_logic;
    AT1_N     : out std_logic;
    TT0_P     : out std_logic;
    TT0_N     : out std_logic;
    TT1_P     : out std_logic;
    TT1_N     : out std_logic;
    
    HMOSI     : in std_logic;
    HMISO     : out std_logic;
    HSCK      : in std_logic;
    HSEL      : in std_logic;
    LA0       : out std_logic_vector (15 downto 0);
    LA1       : out std_logic_vector (15 downto 0);
    LA2       : out std_logic_vector (15 downto 0);
    LA3       : out std_logic_vector (15 downto 0);
    LACK0     : out std_logic;
    LACK1     : out std_logic;
    LACK2     : out std_logic;
    LACK3     : out std_logic;
    EVNT      : out std_logic;
    LED1      : out std_logic;
    LED2      : out std_logic;
    LED3      : out std_logic;
    LED4      : out std_logic;
    MGTCLK_P  : in std_logic;
    MGTCLK_N  : in std_logic;
    GBT_RX_P  : in std_logic;
    GBT_RX_N  : in std_logic;
    GBT_TX_P  : out std_logic;
    GBT_TX_N  : out std_logic;
    FSEL      : out std_logic;
    FMOSI     : out std_logic;
    FMISO     : in std_logic

  );
end PM12;
architecture RTL of PM12 is

  type data_vector is array (0 to 11) of std_logic_vector (32 downto 0);
  type trig_ampl is array (0 to 11) of std_logic_vector(10 downto 0);

  signal RESET, lock320, lock300_1, lock300_2, lock300_3, sreset, rsti, SPI_CS, spi_rd, spi_rden, spi_lock320, spi_lock320_0, hspi_lock320, hspi_lock320_0, cnt_rst, cnt_rd, spi_wr_rdy, spi_wr0, spi_wr1, spi_wr2, spi_wr_req                                                                                : std_logic := '0';
  signal spi_lock_1, spi_lock0_1, spi_lock_2, spi_lock0_2, spi_lock_3, spi_lock0_3, rd_lock_spi, rd_lock_hspi, rd_lock, dcs_irq                                                                                                                                                                               : std_logic;
  signal rstcount                                                                                                                                                                                                                                                                                             : std_logic_vector (3 downto 0);
  signal irq_cnt                                                                                                                                                                                                                                                                                              : std_logic_vector (1 downto 0);
  signal hspi_rden, hcnt_rd, hspi_wr_rdy, hspi_rd, hspi_wr0, hspi_wr1, hspi_wr2, hspi_wr_req, hspibuf_wr, spibuf_wr, hspibuf_rd, spibuf_rd, hspi_na, spi_na, hspi_h                                                                                                                                           : std_logic;
  signal hspibuf_wr0, spibuf_wr0, hspibuf_rd0, spibuf_rd0, hspibuf_wr1, spibuf_wr1, hspibuf_rd1, spibuf_rd1, hspibuf_wr2, spibuf_wr2, hspibuf_rd2, spibuf_rd2                                                                                                                                                 : std_logic;
  signal sbuf_wrena, hbuf_wrena, sbuf_rdena, hbuf_rdena, sbuf_ena, hbuf_ena, hbuf_req, buf_lock, buf_lock0, buf_lock1, buf_lock2, vect_clr, vect_clr_req                                                                                                                                                      : std_logic;
  signal hspi_buf_out, spi_buf_out                                                                                                                                                                                                                                                                            : std_logic_vector (15 downto 0);
  signal buf_cou                                                                                                                                                                                                                                                                                              : std_logic_vector (7 downto 0);
  signal buf_vector, rd_buf_vector                                                                                                                                                                                                                                                                            : std_logic_vector (59 downto 0);
  signal SPI_DATA, spi_wr_data, HSPI_DATA, hspi_wr_data, hspi_wr_data_l, reg_wr_data, hspi_32l                                                                                                                                                                                                                : std_logic_vector (15 downto 0) := (others => '0');
  signal spi_addr, hspi_addr, reg_wr_addr                                                                                                                                                                                                                                                                     : std_logic_vector (8 downto 0)  := (others => '0');
  signal spi_bit_count, hspi_bit_count                                                                                                                                                                                                                                                                        : std_logic_vector (4 downto 0)  := (others => '0');
  signal gate_time_low, gate_time_high                                                                                                                                                                                                                                                                        : std_logic_vector (7 downto 0)  := (others => '0');
  signal reg32_wr, reg32_wr0, reg32_wr1, reg32_wr2, reg32_rd, reg32_rd0, reg32_rd1, reg32_rd2, reg32_str, reg32_str0, reg32_str1, reg32_str2, str_reg32, reg32_320_wr, reg32_320_wr0, reg32_320_wr1, reg32_320_wr2, reg32_320_str, reg32_320_str0, reg32_320_str1, reg32_320_str2                             : std_logic                      := '0';
  signal CH1A_shift, CH1B_shift, CH1C_shift, CH1D_shift, CH2A_shift, CH2B_shift, CH2C_shift, CH2D_shift, CH3A_shift, CH3B_shift, CH3C_shift, CH3D_shift                                                                                                                                                       : std_logic_vector (11 downto 0) := (others => '0');
  signal CH1_0_zero, CH1_1_zero, CH2_0_zero, CH2_1_zero, CH3_0_zero, CH3_1_zero, CH4_0_zero, CH4_1_zero, CH5_0_zero, CH5_1_zero, CH6_0_zero, CH6_1_zero, CH7_0_zero, CH7_1_zero, CH8_0_zero, CH8_1_zero, CH9_0_zero, CH9_1_zero, CH10_0_zero, CH10_1_zero, CH11_0_zero, CH11_1_zero, CH12_0_zero, CH12_1_zero : std_logic_vector (11 downto 0) := (others => '0');
  signal CH1_0_rg, CH1_1_rg, CH2_0_rg, CH2_1_rg, CH3_0_rg, CH3_1_rg, CH4_0_rg, CH4_1_rg, CH5_0_rg, CH5_1_rg, CH6_0_rg, CH6_1_rg, CH7_0_rg, CH7_1_rg, CH8_0_rg, CH8_1_rg, CH9_0_rg, CH9_1_rg, CH10_0_rg, CH10_1_rg, CH11_0_rg, CH11_1_rg, CH12_0_rg, CH12_1_rg                                                 : std_logic_vector (12 downto 0) := (others => '0');
  signal CH1_0_rc, CH1_1_rc, CH2_0_rc, CH2_1_rc, CH3_0_rc, CH3_1_rc, CH4_0_rc, CH4_1_rc, CH5_0_rc, CH5_1_rc, CH6_0_rc, CH6_1_rc, CH7_0_rc, CH7_1_rc, CH8_0_rc, CH8_1_rc, CH9_0_rc, CH9_1_rc, CH10_0_rc, CH10_1_rc, CH11_0_rc, CH11_1_rc, CH12_0_rc, CH12_1_rc                                                 : std_logic_vector (11 downto 0) := (others => '0');

  signal TDCCLK1, TDCCLK2, TDCCLK3, RDA1, RSA1, RDB1, RSB1, RDC1, RSC1, RDD1, RSD1, RDA2, RSA2, RDB2, RSB2, RDC2, RSC2, RDD2, RSD2, RDA3, RSA3, RDB3, RSB3, RDC3, RSC3, RDD3, RSD3, TDCCLK1L, TDCCLK2L, TDCCLK3L                                                 : std_logic;
  signal CH1, CH2, CH3, CH4, CH5, CH6, CH7, CH8, CH9, CH10, CH11, CH12                                                                                                                                                                                           : std_logic_vector (12 downto 0);
  signal CSTR1, CSTR2, CSTR3, CSTR4, CSTR5, CSTR6, CSTR7, CSTR8, CSTR9, CSTR10, CSTR11, CSTR12, CGE1, CGE2, CGE3, CGE4, CGE5, CGE6, CGE7, CGE8, CGE9, CGE10, CGE11, CGE12, CGE1i, CGE2i, CGE3i, CGE4i, CGE5i, CGE6i, CGE7i, CGE8i, CGE9i, CGE10i, CGE11i, CGE12i : std_logic;
  signal SCKI, MISOI, MOSII, LOCKI, TDCHCLI, TDCHDI, TDCHSI, TDCRSI, TDCALMI                                                                                                                                                                                     : std_logic;
  signal MCLK40, MCLK40_1, MCLK40_0, MCLK40T, mclk1, mclk2, mclk3, MGTCLK                                                                                                                                                                                        : std_logic;
  signal MCLK40_IN1, MCLK40_IN2, MCLK40_IN3                                                                                                                                                                                                                      : std_logic;
  signal AT0, AT1, TT0, TT1                                                                                                                                                                                                                                      : std_logic;
  signal HMOSII, HMISOI, HSCKI, HSELI                                                                                                                                                                                                                            : std_logic;
  signal LA0I, LA1I, LA2I, LA3I                                                                                                                                                                                                                                  : std_logic_vector (15 downto 0) := (others => '0');
  signal LACK0I, LACK1I, LACK2I, LACK3I                                                                                                                                                                                                                          : std_logic;

  signal BC_BITS1, BC_BITS2, BC_BITS3 : std_logic_vector (2 downto 0);
  signal BCOLD1, BCOLD2, BCOLD3       : std_logic_vector (1 downto 0);

  signal BC_PER1, BC_PER2, BC_PER3                                                                                                                                            : std_logic_vector (6 downto 0);
  signal BC_JUMP1, BC_JUMP2, BC_JUMP3, ALM_CLR, almclr10, almclr11, alm_clr1, almclr20, almclr21, alm_clr2, almclr30, almclr31, alm_clr3, IRQI                                : std_logic;
  signal HBC_JUMP1, HBC_JUMP2, HBC_JUMP3, hclr10, hclr11, h_clr1, hclr20, hclr21, h_clr2, hclr30, hclr31, h_clr3, Hs_rd, HGBTRXerr, hstat_clr, hstat_clr0, hstat_clr1, Hs_clr : std_logic;

  signal TDC_COU1, TDC_COU2, TDC_COU3 : std_logic_vector (3 downto 0) := (others => '0');

  signal TDC1A, TDC1B, TDC1C, TDC1D, TDC2A, TDC2B, TDC2C, TDC2D, TDC3A, TDC3B, TDC3C, TDC3D : std_logic_vector (11 downto 0);

  signal CH_TIME_T : trig_time;
  --signal Trig_on0, Trig_onA0 : STD_LOGIC;
  signal GBT_TX_D, GBT_RX_D : std_logic_vector (79 downto 0);

  signal TDC1A_raw, TDC1B_raw, TDC1C_raw, TDC1D_raw, TDC2A_raw, TDC2B_raw, TDC2C_raw, TDC2D_raw, TDC3A_raw, TDC3B_raw, TDC3C_raw, TDC3D_raw : std_logic_vector (12 downto 0);

  signal clk300_1, clk300_2, clk300_3, clk600_1, clk600_2, clk600_3, clk600_90_1, clk600_90_2, clk600_90_3, clk320, clkfbin1, clkfbout1, clkfbin2, clkfbout2, clkfbin3, clkfbout3 : std_logic;

  signal BC_STR1, BC_STR11, BC_STR12, BC_STR2, BC_STR21, BC_STR22, BC_STR3, BC_STR31, BC_STR32, C1_EV                                                   : std_logic;
  signal F1A_full, F1B_full, F1C_full, F1D_full, F2A_full, F2B_full, F2C_full, F2D_full, F3A_full, F3B_full, F3C_full, F3D_full, Trig_on0, Trig_onA0    : std_logic;
  signal TDC1A_rdy0, TDC1B_rdy0, TDC1C_rdy0, TDC1D_rdy0, TDC2A_rdy0, TDC2B_rdy0, TDC2C_rdy0, TDC2D_rdy0, TDC3A_rdy0, TDC3B_rdy0, TDC3C_rdy0, TDC3D_rdy0 : std_logic;
  signal mt_cou                                                                                                                                         : std_logic_vector(2 downto 0)  := (others => '0');
  signal BC_cou                                                                                                                                         : std_logic_vector(11 downto 0) := (others => '0');
  signal TR_to                                                                                                                                          : std_logic_vector(5 downto 0)  := (others => '0');

  signal CH_ampl0 : trig_ampl0;

  signal N_chans : std_logic_vector(3 downto 0) := (others => '0');

  signal tt, ta, tto, tao : std_logic_vector (1 downto 0) := (others => '0');

  signal GBT_is_RXD, GBT_is_TXD, RX_CLK, TX_CLK, GBTRX_ready, GBTRX_ready0, GBT_chg, HGBT_chg, GBT_rdy, GBT_rdy0, t100ms, RX_err, RX_err1, RX_err_LED, rxerr0, TXact, RXact, RXLED, TXLED, txled0, rxled0, LNKLED, IsRXData0, GBTRXerr, stat_clr, stat_clr0, stat_clr1 : std_logic;
  signal cou_100ms                                                                                                                                                                                                                                                     : std_logic_vector (21 downto 0);
  signal alm_rst0, alm_rst, chans_block, is_rst                                                                                                                                                                                                                        : std_logic;

  signal chans_ena, chans_ena_r                                                                                                                                                                               : std_logic_vector (11 downto 0) := (others => '0');
  signal CH1_Z0, CH1_Z1, CH2_Z0, CH2_Z1, CH3_Z0, CH3_Z1, CH4_Z0, CH4_Z1, CH5_Z0, CH5_Z1, CH6_Z0, CH6_Z1, CH7_Z0, CH7_Z1, CH8_Z0, CH8_Z1, CH9_Z0, CH9_Z1, CH10_Z0, CH10_Z1, CH11_Z0, CH11_Z1, CH12_Z0, CH12_Z1 : std_logic_vector (15 downto 0);

  signal N1_chans, N2_chans : std_logic_vector (2 downto 0);
  signal TT_mode            : std_logic;

  signal ampl_sat                                                                                                                                                            : std_logic_vector (11 downto 0) := (others => '0');
  signal ampl_low                                                                                                                                                            : std_logic_vector (3 downto 0)  := (others => '0');
  signal Event_in, DATA_rd, DATA_rdy, inp_cou, CH_trig, CH_triga, CH_do, Z_alarm, trig_bgnd, cnt_trig, trig_dis, ch_trig_outtn                                               : std_logic_vector (11 downto 0) := (others => '0');
  signal inp_event, EV_ID_wr, EV_ID_rd, EV_ID_empty, Event_ready, Event_ready_0, Event_free, wr_out_id, New_BCID, DATA80_rd, DATA_empty, FIFO_dis, wr_nch, ev_tout, ev_tout0 : std_logic;
  signal ev_tout_cnt                                                                                                                                                         : std_logic_vector (7 downto 0);

  signal CH_N0, CH_N1, CH_N0_0, CH_N1_0, CH_NUM                                                                                                                                     : std_logic_vector (3 downto 0);
  signal CH_NUM1, CH_NUM2                                                                                                                                                           : std_logic_vector (2 downto 0);
  signal WRDS_NUM                                                                                                                                                                   : std_logic_vector (2 downto 0);
  signal Orbit_ID, hspid_w32, hspid_r32, tstamp, hspib_32, mcu_tstamp                                                                                                               : std_logic_vector (31 downto 0);
  signal xadc_r, xadc_out                                                                                                                                                           : std_logic_vector (15 downto 0);
  signal xadc_a                                                                                                                                                                     : std_logic_vector (6 downto 0);
  signal EV_ID_in, EV_ID_out                                                                                                                                                        : std_logic_vector (55 downto 0);
  signal EV_DATA80, DATA80_in, data_word                                                                                                                                            : std_logic_vector (79 downto 0);
  signal is_data, is_header                                                                                                                                                         : std_logic;
  signal WR_fifo_out, wr_hspi32, rd_hspi32, flsh_sel, TCM_req, TCM_reqh, TCM_req0, TCM_req1, TCM_req2, fl_rst, rd_xadc, xadc_en, xadc_rdy, gs0_0, gs1_0, gs0_1, gs1_1, rdo_sel, fdd : std_logic := '0';

  signal DATA_out          : data_vector;
  signal ev_out_cou        : std_logic_vector (3 downto 0);
  signal cnt_out, hcnt_out : std_logic_vector (15 downto 0);

  signal psen1, psincdec1, jumpa1, flock1, fdone1, psen2, psincdec2, jumpa2, flock2, fdone2, psen3, psincdec3, jumpa3, flock3, fdone3, all_locked : std_logic;
  signal pshift1, pshift2, pshift3                                                                                                                : std_logic_vector (5 downto 0);

  signal rx_phase_status : std_logic_vector(3 downto 0);

  signal hyst_md                                                                                      : std_logic_vector(15 downto 0);
  signal start_hyst, h_busy, wr_hyst_a, rd_hyst_d, hysta_sel, hystd_sel, hyst_stp, hyst_rst, hyst_clr : std_logic;
  signal cnt_md                                                                                       : std_logic := '0';
  signal hyst_data                                                                                    : hyst_vector;
  signal hyst_a, hyst_t                                                                               : std_logic_vector(11 downto 0);
  signal hyst_addr                                                                                    : std_logic_vector(16 downto 0);
  signal hyst_r_data                                                                                  : std_logic_vector(31 downto 0);
  component PLL320
    port
    (
      mclk_in : in std_logic;
      RESET   : in std_logic;
      locked  : out std_logic;
      CLK320  : out std_logic;
      CLK40   : out std_logic);
  end component;

  component CLK600_pll
    port
    (
      CLK_IN    : in std_logic;
      RESET     : in std_logic;
      CLKFB_IN  : in std_logic;
      locked    : out std_logic;
      psclk     : in std_logic;
      psen      : in std_logic;
      psincdec  : in std_logic;
      psdone    : out std_logic;
      CLK600    : out std_logic;
      CLK600_90 : out std_logic;
      CLK300    : out std_logic;
      CLKFB_OUT : out std_logic);
  end component;

  component pin_capt
    port
    (
      pin_in    : in std_logic;
      pin_out   : out std_logic;
      clk600    : in std_logic;
      clk600_90 : in std_logic;
      clk300    : in std_logic;
      str       : out std_logic;
      ptime     : out std_logic_vector (2 downto 0));
  end component;

  component TDCCHAN is
    port
    (
      pin_in    : in std_logic;
      pin_out   : out std_logic;
      clk300    : in std_logic;
      clk600    : in std_logic;
      clk600_90 : in std_logic;
      reset     : in std_logic;
      tdcclk    : in std_logic;
      rstr      : in std_logic;
      rdata     : in std_logic;
      tdc_count : in std_logic_vector (3 downto 0);
      bc_time   : in std_logic_vector (6 downto 0);
      tdc_out   : out std_logic_vector (11 downto 0);
      tdc_rdy   : out std_logic;
      --             fifo_full : out STD_LOGIC;
      tdc_raw      : out std_logic_vector (12 downto 0);
      tdc_raw_lock : in std_logic
    );
  end component;

  component Channel is
    port
    (
      CGE        : in std_logic;
      clk320     : in std_logic;
      reset      : in std_logic;
      tdc_rdy_in : in std_logic;
      mt_cou     : in std_logic_vector (2 downto 0);
      bc_cou     : in std_logic_vector (5 downto 0);
      TR_bc      : in std_logic_vector (5 downto 0);
      TDC        : in std_logic_vector (11 downto 0);
      --              TDC_full : in STD_LOGIC;
      CSTR           : in std_logic;
      CH             : in std_logic_vector(12 downto 0);
      CH_shift       : in std_logic_vector (11 downto 0);
      gate_time_low  : in std_logic_vector (7 downto 0);
      FIFO_dis       : in std_logic;
      gate_time_high : in std_logic_vector (7 downto 0);
      Ampl_sat       : in std_logic_vector (11 downto 0);
      ampl_low       : in std_logic_vector (3 downto 0);
      CH0_zero       : out std_logic_vector (11 downto 0);
      CH1_zero       : out std_logic_vector (11 downto 0);
      CH_trig_outt   : out std_logic;
      CH_trig_outa   : out std_logic;
      CH_trig_bgnd   : out std_logic;
      CH_TIME        : out std_logic_vector (9 downto 0);
      CH_ampl        : out std_logic_vector (12 downto 0);
      DATA_out       : out std_logic_vector (32 downto 0);
      DATA_ready     : out std_logic;
      DATA_rd        : in std_logic;
      Event_in       : out std_logic;
      Z0_cal         : out std_logic_vector (15 downto 0);
      Z1_cal         : out std_logic_vector (15 downto 0);
      Z_alarm        : out std_logic;
      spi_lock       : in std_logic;
      R0_cal         : out std_logic_vector (12 downto 0);
      R1_cal         : out std_logic_vector (12 downto 0);
      R0_corr        : in std_logic_vector (11 downto 0);
      R1_corr        : in std_logic_vector (11 downto 0);
      pulse_in       : out std_logic;
      chan_ena       : in std_logic;
      trig_dis       : in std_logic;
      fdd            : in std_logic;
      CH_trig_int    : in std_logic;
      CH_trig_outtn  : out std_logic
    );

  end component;

  component EVENTID_FIFO
    port
    (
      clk   : in std_logic;
      srst  : in std_logic;
      din   : in std_logic_vector(55 downto 0);
      wr_en : in std_logic;
      rd_en : in std_logic;
      dout  : out std_logic_vector(55 downto 0);
      full  : out std_logic;
      empty : out std_logic);
  end component;
  -- ###############################################
  -- #########  GBT Readout ########################
  -- ###############################################
  signal readout_status    : readout_status_t;
  signal readout_control   : readout_control_t;
  signal Data_from_FITrd   : std_logic_vector(GBT_data_word_bitdepth - 1 downto 0);
  signal IsData_from_FITrd : std_logic;

  signal RxData_rxclk_from_GBT   : std_logic_vector(GBT_data_word_bitdepth - 1 downto 0);
  signal IsRxData_rxclk_from_GBT : std_logic;

  signal PM_data_toreadout : board_data_type;

  signal ipbus_control_reg : ctrl_reg_t;
  signal ipbus_status_reg  : stat_reg_t;

  signal gbt_global_status    : std_logic_vector(3 downto 0);
  signal err_report_fifo_rden : std_logic;
  signal readout_err_rden     : std_logic;

  component FIT_GBT_project is
    generic
    (
      IS_SIMULATION : integer := 0
    );

    port
    (
      RESET_I          : in std_logic;
      SysClk_I         : in std_logic; -- 320MHz system clock
      DataClk_I        : in std_logic; -- 40MHz data clock
      MgtRefClk_I      : in std_logic; -- 200MHz ref clock
      RxDataClk_I      : in std_logic; -- 40MHz data clock in RX domain
      GBT_RxFrameClk_O : out std_logic; --Rx GBT frame clk 40MHz
      FSM_Clocks_O     : out rdclocks_t;

      IPbusClk_I             : in std_logic; -- IPbus clock for error fifo read
      err_report_fifo_rden_i : in std_logic; -- IPbus error report fifo read enable

      Board_data_I       : in board_data_type; --PM or TCM data
      Control_register_I : in readout_control_t;
      errors_rden_I      : in std_logic; -- status register EA (errors) was read

      MGT_RX_P_I    : in std_logic;
      MGT_RX_N_I    : in std_logic;
      MGT_TX_P_O    : out std_logic;
      MGT_TX_N_O    : out std_logic;
      MGT_TX_dsbl_O : out std_logic;

      -- GBT data to/from FIT readout 
      RxData_rxclk_to_FITrd_I   : in std_logic_vector(GBT_data_word_bitdepth - 1 downto 0);
      IsRxData_rxclk_to_FITrd_I : in std_logic;
      Data_from_FITrd_O         : out std_logic_vector(GBT_data_word_bitdepth - 1 downto 0);
      IsData_from_FITrd_O       : out std_logic;

      -- GBT data to/from GBT project
      Data_to_GBT_I             : in std_logic_vector(GBT_data_word_bitdepth - 1 downto 0);
      IsData_to_GBT_I           : in std_logic;
      RxData_rxclk_from_GBT_O   : out std_logic_vector(GBT_data_word_bitdepth - 1 downto 0);
      IsRxData_rxclk_from_GBT_O : out std_logic;
      -- FIT readour status, including BCOR_ID to PM/TCM
      readout_status_o : out readout_status_t

    );
  end component;
  -- ###############################################
  -- ###############################################
  -- ###############################################
  component counters
    port
    (
      clk    : in std_logic;
      evnt   : in std_logic_vector (11 downto 0);
      trig   : in std_logic_vector (11 downto 0);
      reset  : in std_logic;
      dout   : out std_logic_vector (15 downto 0);
      hdout  : out std_logic_vector (15 downto 0);
      raddr  : in std_logic_vector (5 downto 0);
      hraddr : in std_logic_vector (4 downto 0);
      hl     : in std_logic;
      rd_en  : in std_logic;
      hrd_en : in std_logic
    );
  end component;

  component trigger
    port
    (
      clk320    : in std_logic;
      mt_cou    : in std_logic_vector (2 downto 0);
      CH_trigt  : in std_logic_vector (11 downto 0);
      CH_triga  : in std_logic_vector (11 downto 0);
      CH_trigb  : in std_logic_vector (11 downto 0);
      CH_TIME_T : in trig_time;
      CH_ampl0  : in trig_ampl0;
      tcm_req   : in std_logic;
      tt        : out std_logic_vector (1 downto 0);
      ta        : out std_logic_vector (1 downto 0)
    );
  end component;

  component Xmega_buf
    port
    (
      clka  : in std_logic;
      ena   : in std_logic;
      wea   : in std_logic_vector(0 downto 0);
      addra : in std_logic_vector(5 downto 0);
      dina  : in std_logic_vector(15 downto 0);
      douta : out std_logic_vector(15 downto 0);
      clkb  : in std_logic;
      enb   : in std_logic;
      web   : in std_logic_vector(0 downto 0);
      addrb : in std_logic_vector(5 downto 0);
      dinb  : in std_logic_vector(15 downto 0);
      doutb : out std_logic_vector(15 downto 0)
    );
  end component;

  component FLASH
    generic
    (
      clk_freq : integer
    );
    port
    (
      rst         : in std_logic;
      clk         : in std_logic;
      data_in     : in std_logic_vector(31 downto 0);
      data_out    : out std_logic_vector(31 downto 0);
      A           : in std_logic_vector(1 downto 0);
      wr_flshreg  : in std_logic;
      rd_flshreg  : in std_logic;
      flshreg_sel : in std_logic;
      FSEL        : out std_logic;
      FMOSI       : out std_logic;
      FMISO       : in std_logic
    );
  end component;

  component SENSOR
    port
    (
      di_in       : in std_logic_vector(15 downto 0);
      daddr_in    : in std_logic_vector(6 downto 0);
      den_in      : in std_logic;
      dwe_in      : in std_logic;
      drdy_out    : out std_logic;
      do_out      : out std_logic_vector(15 downto 0);
      dclk_in     : in std_logic;
      reset_in    : in std_logic;
      vp_in       : in std_logic;
      vn_in       : in std_logic;
      channel_out : out std_logic_vector(4 downto 0);
      eoc_out     : out std_logic;
      alarm_out   : out std_logic;
      eos_out     : out std_logic;
      busy_out    : out std_logic
    );
  end component;

  component autophase
    port
    (
      clk      : in std_logic;
      lock     : in std_logic;
      jump     : in std_logic;
      psen     : out std_logic;
      psincdec : out std_logic;
      done     : out std_logic;
      shift    : out std_logic_vector (5 downto 0)
    );
  end component;

  component hyst
    port
    (
      clk320        : in std_logic;
      hyst_inp_data : in hyst_vector;
      hyst_a        : in std_logic_vector(11 downto 0);
      hyst_t        : in std_logic_vector(11 downto 0);
      hyst_st       : in std_logic;
      cnt_clr       : in std_logic;
      busy          : out std_logic;
      hyst_addr_i   : in std_logic_vector(16 downto 0);
      hyst_addr_o   : out std_logic_vector(16 downto 0);
      wr_addr       : in std_logic;
      hyst_data_o   : out std_logic_vector(31 downto 0);
      n_addr        : in std_logic;
      lock320       : in std_logic;
      stp           : out std_logic
    );
  end component;

  -- attribute mark_debug              : string;
  -- attribute mark_debug of rd_hspi32     : signal is "true";
  -- attribute mark_debug of hspib_32     : signal is "true";
  -- attribute mark_debug of hspi_addr     : signal is "true";
  -- attribute mark_debug of err_report_fifo_rden     : signal is "true";
  -- attribute mark_debug of readout_err_rden     : signal is "true";

begin

  TCLK1 : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port map
    (I => TDCCLK1_P, IB => TDCCLK1_N, O => TDCCLK1L);

  TCLKB1 : BUFR
  generic
  map (BUFR_DIVIDE => "BYPASS")
  port
  map (O => TDCCLK1, CE => '1', CLR => '0', I => TDCCLK1L);

  TCLK2 : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => TDCCLK2_P, IB => TDCCLK2_N, O => TDCCLK2L);

  TCLKB2 : BUFR
  generic
  map (BUFR_DIVIDE => "BYPASS")
  port
  map (O => TDCCLK2, CE => '1', CLR => '0', I => TDCCLK2L);

  TCLK3 : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => TDCCLK3_P, IB => TDCCLK3_N, O => TDCCLK3L);

  TCLKB3 : BUFR
  generic
  map (BUFR_DIVIDE => "BYPASS")
  port
  map (O => TDCCLK3, CE => '1', CLR => '0', I => TDCCLK3L);
  RDA1_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RDA1_P, IB => RDA1_N, O => RDA1);
  RSA1_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RSA1_P, IB => RSA1_N, O => RSA1);
  RDB1_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RDB1_P, IB => RDB1_N, O => RDB1);
  RSB1_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RSB1_P, IB => RSB1_N, O => RSB1);
  RDC1_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RDC1_P, IB => RDC1_N, O => RDC1);
  RSC1_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RSC1_P, IB => RSC1_N, O => RSC1);
  RDD1_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RDD1_P, IB => RDD1_N, O => RDD1);
  RSD1_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RSD1_P, IB => RSD1_N, O => RSD1);

  RDA2_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RDA2_P, IB => RDA2_N, O => RDA2);
  RSA2_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RSA2_P, IB => RSA2_N, O => RSA2);
  RDB2_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RDB2_P, IB => RDB2_N, O => RDB2);
  RSB2_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RSB2_P, IB => RSB2_N, O => RSB2);
  RDC2_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RDC2_P, IB => RDC2_N, O => RDC2);
  RSC2_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RSC2_P, IB => RSC2_N, O => RSC2);
  RDD2_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RDD2_P, IB => RDD2_N, O => RDD2);
  RSD2_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RSD2_P, IB => RSD2_N, O => RSD2);

  RDA3_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RDA3_P, IB => RDA3_N, O => RDA3);
  RSA3_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RSA3_P, IB => RSA3_N, O => RSA3);
  RDB3_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RDB3_P, IB => RDB3_N, O => RDB3);
  RSB3_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RSB3_P, IB => RSB3_N, O => RSB3);
  RDC3_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RDC3_P, IB => RDC3_N, O => RDC3);
  RSC3_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RSC3_P, IB => RSC3_N, O => RSC3);
  RDD3_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RDD3_P, IB => RDD3_N, O => RDD3);
  RSD3_B : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => RSD3_P, IB => RSD3_N, O => RSD3);
  ADCIN : for i in 0 to 12 generate
    ADC1 : IBUF
    port
    map (O => CH1(i), I => DI1(i));
    ADC2 : IBUF
    port
    map (O => CH2(i), I => DI2(i));
    ADC3 : IBUF
    port
    map (O => CH3(i), I => DI3(i));
    ADC4 : IBUF
    port
    map (O => CH4(i), I => DI4(i));
    ADC5 : IBUF
    port
    map (O => CH5(i), I => DI5(i));
    ADC6 : IBUF
    port
    map (O => CH6(i), I => DI6(i));
    ADC7 : IBUF
    port
    map (O => CH7(i), I => DI7(i));
    ADC8 : IBUF
    port
    map (O => CH8(i), I => DI8(i));
    ADC9 : IBUF
    port
    map (O => CH9(i), I => DI9(i));
    ADC10 : IBUF
    port
    map (O => CH10(i), I => DI10(i));
    ADC11 : IBUF
    port
    map (O => CH11(i), I => DI11(i));
    ADC12 : IBUF
    port
    map (O => CH12(i), I => DI12(i));
  end generate;

  iN1 : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => INA1_P, IB => INA1_N, O => CGE1i);
  iN2 : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => INB1_P, IB => INB1_N, O => CGE2i);
  iN3 : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => INC1_P, IB => INC1_N, O => CGE3i);
  iN4 : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => IND1_P, IB => IND1_N, O => CGE4i);
  iN5 : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => INA2_P, IB => INA2_N, O => CGE5i);
  iN6 : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => INB2_P, IB => INB2_N, O => CGE6i);
  iN7 : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => INC2_P, IB => INC2_N, O => CGE7i);
  iN8 : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => IND2_P, IB => IND2_N, O => CGE8i);
  iN9 : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => INA3_P, IB => INA3_N, O => CGE9i);
  iN10 : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => INB3_P, IB => INB3_N, O => CGE10i);
  iN11 : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => INC3_P, IB => INC3_N, O => CGE11i);
  iN12 : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => IND3_P, IB => IND3_N, O => CGE12i);
  iSTR1 : IBUF
  port
  map (O => CSTR1, I => STR1);
  iSTR2 : IBUF
  port
  map (O => CSTR2, I => STR2);
  iSTR3 : IBUF
  port
  map (O => CSTR3, I => STR3);
  iSTR4 : IBUF
  port
  map (O => CSTR4, I => STR4);
  iSTR5 : IBUF
  port
  map (O => CSTR5, I => STR5);
  iSTR6 : IBUF
  port
  map (O => CSTR6, I => STR6);
  iSTR7 : IBUF
  port
  map (O => CSTR7, I => STR7);
  iSTR8 : IBUF
  port
  map (O => CSTR8, I => STR8);
  iSTR9 : IBUF
  port
  map (O => CSTR9, I => STR9);
  iSTR10 : IBUF
  port
  map (O => CSTR10, I => STR10);
  iSTR11 : IBUF
  port
  map (O => CSTR11, I => STR11);
  iSTR12 : IBUF
  port
  map (O => CSTR12, I => STR12);

  iSCK : IBUF
  port
  map (O => SCKI, I => SCK);
  iMISO : OBUFT
  port
  map (I => MISOI, O => MISO, T => spi_rden);
  iMOSI : IBUF
  port
  map (O => MOSII, I => MOSI);
  iCS : IBUF
  port
  map (O => SPI_CS, I => CS);
  iRST : IBUF
  port
  map (O => rsti, I => RST);

  iMCLK1 : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => MCLK1_P, IB => MCLK1_N, O => MCLK1);

  iMCLK2 : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => MCLK2_P, IB => MCLK2_N, O => MCLK2);

  iMCLK3 : IBUFDS
  generic
  map (DIFF_TERM => TRUE, IBUF_LOW_PWR => FALSE, IOSTANDARD => "LVDS")
  port
  map (I => MCLK3_P, IB => MCLK3_N, O => MCLK3);

  iAT0 : OBUFDS
  generic
  map (SLEW => "FAST", IOSTANDARD => "LVDS") port
  map (I => AT0, OB => AT0_N, O => AT0_P);
  iAT1 : OBUFDS
  generic
  map (SLEW => "FAST", IOSTANDARD => "LVDS") port
  map (I => AT1, OB => AT1_N, O => AT1_P);
  iTT0 : OBUFDS
  generic
  map (SLEW => "FAST", IOSTANDARD => "LVDS") port
  map (I => TT0, OB => TT0_N, O => TT0_P);
  iTT1 : OBUFDS
  generic
  map (SLEW => "FAST", IOSTANDARD => "LVDS") port
  map (I => TT1, OB => TT1_N, O => TT1_P);

  iHMOSI : IBUF
  port
  map (O => HMOSII, I => HMOSI);
  iHSCK : IBUF
  port
  map (O => HSCKI, I => HSCK);
  iHSEL : IBUF
  port
  map (O => HSELI, I => HSEL);
  iHMISO : OBUFT
  port
  map (O => HMISO, I => HMISOI, T => hspi_rden);

  ILA : for i in 0 to 15 generate
    ILA0 : OBUF
    port
    map (O => LA0(i), I => LA0I(i));
    ILA1 : OBUF
    port
    map (O => LA1(i), I => LA1I(i));
    ILA2 : OBUF
    port
    map (O => LA2(i), I => LA2I(i));
    ILA3 : OBUF
    port
    map (O => LA3(i), I => LA3I(i));
  end generate;

  ILACK0 : OBUF
  port
  map (O => LACK0, I => LACK0I);
  ILACK1 : OBUF
  port
  map (O => LACK1, I => LACK1I);
  ILACK2 : OBUF
  port
  map (O => LACK2, I => LACK2I);
  ILACK3 : OBUF
  port
  map (O => LACK3, I => LACK3I);

  ILED1 : OBUF
  port
  map (O => LED1, I => TXLED);
  ILED2 : OBUF
  port
  map (O => LED2, I => RXLED);
  ILED3 : OBUF
  port
  map (O => LED3, I => LNKLED);
  ILED4 : OBUF
  port
  map (O => LED4, I => RX_err_LED);
  IRQ1 : OBUF
  port
  map (O => IRQ, I => IRQI);

  IEVNT : OBUF
  port
  map (O => EVNT, I => '0');

  IMGTCLK1 : IBUFDS_GTE2
  port
  map (O => MGTCLK, I => MGTCLK_P, IB => MGTCLK_N, CEB => '0');

  fl_upg : FLASH generic
  map (clk_freq => 40000)
  port
  map (rst => fl_rst, clk => TX_CLK, data_in => hspid_w32, data_out => hspid_r32, A => hspi_addr(1 downto 0), wr_flshreg => wr_hspi32, rd_flshreg => str_reg32, flshreg_sel => flsh_sel, FSEL => FSEL, FMOSI => FMOSI, FMISO => FMISO);
  IRQI <= BC_JUMP1 or BC_JUMP2 or BC_JUMP3 or GBTRXerr or GBT_chg or dcs_irq when (irq_cnt = "11") else
    '0';

  at0 <= tao(0);
  at1 <= tao(1);
  tt0 <= tto(0);
  tt1 <= tto(1);

  -- #################################################################################################
  -- #################   FIT GBT Readout    ##########################################################
  -- #################################################################################################
  --GBT1:  GBT_TX_RX port map (
  --            RESET =>RESET, 
  --            MgtRefClk => MGTCLK, 
  --            MGT_RX_P =>GBT_RX_P,
  --            MGT_RX_N =>GBT_RX_N,  
  --            MGT_TX_P =>GBT_TX_P, 
  --            MGT_TX_N =>GBT_TX_N, 
  --            TXDataClk =>TX_CLK, 
  --            TXData => GBT_TX_D, 
  --            TXData_SC=>"0000", 
  --            IsTXData =>GBT_is_TXD, 
  --            RXDataClk => RX_CLK, 
  --            RXData =>GBT_RX_D, 
  --            RXData_SC =>open, 
  --            IsRXData => GBT_is_RXD, 
  --            RX_ready=>GBTRX_ready, 
  --            RX_errors=> RX_err
  --        );

  -- FIT GBT project =====================================
  FitGbtPrg : FIT_GBT_project
  generic
  map(
  IS_SIMULATION => 0
  )

  port
  map(
  RESET_I          => sreset,
  SysClk_I         => clk320,
  DataClk_I        => TX_CLK,
  MgtRefClk_I      => MGTCLK,
  RxDataClk_I      => RX_CLK, -- 40MHz data clock in RX domain (loop back)
  GBT_RxFrameClk_O => RX_CLK,
  FSM_Clocks_O     => open,

  IPbusClk_I             => TX_CLK,
  err_report_fifo_rden_i => err_report_fifo_rden,

  Board_data_I       => PM_data_toreadout,
  Control_register_I => readout_control,
  errors_rden_I      => readout_err_rden,

  MGT_RX_P_I    => GBT_RX_P,
  MGT_RX_N_I    => GBT_RX_N,
  MGT_TX_P_O    => GBT_TX_P,
  MGT_TX_N_O    => GBT_TX_N,
  MGT_TX_dsbl_O => open,

  RxData_rxclk_to_FITrd_I   => RxData_rxclk_from_GBT, --loop back data
  IsRxData_rxclk_to_FITrd_I => IsRxData_rxclk_from_GBT, --loop back data
  Data_from_FITrd_O         => Data_from_FITrd,
  IsData_from_FITrd_O       => IsData_from_FITrd,
  Data_to_GBT_I             => Data_from_FITrd, --loop back data
  IsData_to_GBT_I           => IsData_from_FITrd, --loop back data

  RxData_rxclk_from_GBT_O   => RxData_rxclk_from_GBT,
  IsRxData_rxclk_from_GBT_O => IsRxData_rxclk_from_GBT,

  readout_status_o => readout_status
  );
  -- =====================================================

  GBTRX_ready <= readout_status.GBT_status.gbtRx_Ready;
  GBT_is_RXD  <= IsRxData_rxclk_from_GBT;
  RX_err      <= readout_status.GBT_status.gbtRx_ErrorDet;

  --PM_data_toreadout.is_header  <=  GBT_is_TXD;
  --PM_data_toreadout.is_data    <=  GBT_is_TXD;
  --PM_data_toreadout.is_packet  <=  GBT_is_TXD;
  --PM_data_toreadout.data_word  <=  GBT_TX_D;
  readout_control  <= func_CNTRREG_getcntrreg(ipbus_control_reg);
  ipbus_status_reg <= func_STATREG_getaddrreg(readout_status);

  gbt_global_status(0) <= readout_status.Rx_Phase_error;
  gbt_global_status(1) <= '1' when readout_status.BCIDsync_Mode = mode_LOST else
  '0';
  --gbt_global_status(2) <=  '1' when readout_status.hits_rd_counter_selector.hits_skipped /= x"0000_0000" else '0';
  gbt_global_status(3) <= '0';

  process (clk320)
  begin
    if (clk320'event and clk320 = '1') then
      if (readout_status.fsm_errors = x"00") then
        gbt_global_status(2) <= '0';
      else
        gbt_global_status(2) <= '1';
      end if;
      if (cnt_md = '0') then
        cnt_trig <= CH_trig;
      else
        cnt_trig <= CH_triga;
      end if;

    end if;

  end process;
  --gbt_global_status <=  x"0";

  -- #################################################################################################
  -- #################################################################################################

  LNKLED     <= not GBTRX_ready;
  RX_err_LED <= rxerr0 or (not GBTRX_ready);
  TXLED      <= txled0 or (not GBTRX_ready);
  RXLED      <= rxled0 or (not GBTRX_ready);
  process (TX_CLK)
  begin
    if (TX_CLK'event and TX_CLK = '1') then

      if (xadc_rdy = '1') then
        xadc_r <= xadc_out;
      end if;

      fl_rst <= sreset;

      GBT_is_TXD   <= IsData_from_FITrd;
      IsRXData0    <= GBT_is_RXD;
      GBTRX_ready0 <= GBTRX_ready;

      stat_clr0  <= ALM_CLR;
      stat_clr1  <= stat_clr0;
      stat_clr   <= stat_clr1;
      hstat_clr0 <= Hs_rd;
      hstat_clr1 <= hstat_clr0;
      hstat_clr  <= hstat_clr1;
      if (stat_clr1 = '1') and (stat_clr = '0') then
        irq_cnt <= "00";
      else
        if (irq_cnt /= "11") then
          irq_cnt <= irq_cnt + 1;
        end if;
      end if;

      if (GBTRX_ready /= GBTRX_ready0) then
        GBT_chg  <= '1';
        HGBT_chg <= '1';
      else
        if (stat_clr1 = '1') and (stat_clr = '0') then
          GBT_chg <= '0';
        end if;
        if (hstat_clr1 = '1') and (hstat_clr = '0') then
          HGBT_chg <= '0';
        end if;
      end if;

      if (GBTRX_ready = '1') and (GBT_rdy = '1') and (RX_err = '1') then
        GBTRXerr  <= '1';
        HGBTRXerr <= '1';
      else
        if (stat_clr1 = '1') and (stat_clr = '0') then
          GBTRXerr <= '0';
        end if;
        if (hstat_clr1 = '1') and (hstat_clr = '0') then
          HGBTRXerr <= '0';
        end if;
      end if;

      if GBTRX_ready = '0' then
        GBT_rdy0 <= '0';
        GBT_rdy  <= '0';
      else
        if (t100ms = '1') then
          GBT_rdy0 <= '1';
          if (GBT_rdy0 = '1') then
            GBT_rdy <= '1';
          end if;
        end if;
      end if;
      if t100ms = '0' then
        cou_100ms <= cou_100ms + 1;
        if RX_err = '1' then
          RX_err1 <= '1';
        end if;
        if GBT_is_TXD = '1' then
          TXact <= '1';
        end if;
        if IsRXData0 = '1' then
          RXact <= '1';
        end if;
      else
        cou_100ms <= "00" & x"00000";
        RX_err1   <= '0';
        TXact     <= '0';
        RXact     <= '0';
        if (RX_err = '1') or (RX_err1 = '1') then
          RXerr0 <= '0';
        else
          RXerr0 <= '1';
        end if;
        if (GBT_is_TXD = '1') or (TXact = '1') then
          txled0 <= '0';
        else
          txled0 <= '1';
        end if;
        if (IsRXData0 = '1') or (RXact = '1') then
          rxled0 <= '0';
        else
          rxled0 <= '1';
        end if;
      end if;
    end if;
  end process;

  t100ms <= '1' when cou_100ms = "11" & x"D08FF" else
    '0';

  MCLKB1 : BUFR
  generic
  map (
  BUFR_DIVIDE => "BYPASS"
  )
  port
  map (
  O   => MCLK40,
  CE  => '1',
  CLR => '0',
  I   => MCLK40_IN1
  );

  process (MCLK40)
  begin
    if (MCLK40'event and MCLK40 = '1') then
      MCLK40T <= not MCLK40T;
    end if;
  end process;

  af1 : autophase port
  map(clk => clk300_1, lock => flock1, jump => jumpa1, psen => psen1, psincdec => psincdec1, done => fdone1, shift => pshift1);
  PLL1 : CLK600_pll port
  map(CLK_IN => MCLK40_IN1, RESET => RESET, CLKFB_IN => clkfbin1, locked => flock1, psclk => clk300_1, psen => psen1, psincdec => psincdec1, psdone => open, CLK600 => clk600_1, CLK600_90 => CLK600_90_1, CLK300 => clk300_1, CLKFB_OUT => clkfbout1);
  FBBUF1 : BUFH port
  map(O => clkfbin1, I => clkfbout1);
  af2 : autophase port
  map(clk => clk300_2, lock => flock2, jump => jumpa2, psen => psen2, psincdec => psincdec2, done => fdone2, shift => pshift2);
  PLL2 : CLK600_pll port
  map(CLK_IN => MCLK40_IN2, RESET => RESET, CLKFB_IN => clkfbin2, locked => flock2, psclk => clk300_2, psen => psen2, psincdec => psincdec2, psdone => open, CLK600 => clk600_2, CLK600_90 => CLK600_90_2, CLK300 => clk300_2, CLKFB_OUT => clkfbout2);
  FBBUF2 : BUFH port
  map(O => clkfbin2, I => clkfbout2);
  af3 : autophase port
  map(clk => clk300_3, lock => flock3, jump => jumpa3, psen => psen3, psincdec => psincdec3, done => fdone3, shift => pshift3);
  PLL3 : CLK600_pll port
  map(CLK_IN => MCLK40_IN3, RESET => RESET, CLKFB_IN => clkfbin3, locked => flock3, psclk => clk300_3, psen => psen3, psincdec => psincdec3, psdone => open, CLK600 => clk600_3, CLK600_90 => CLK600_90_3, CLK300 => clk300_3, CLKFB_OUT => clkfbout3);
  FBBUF3 : BUFH port
  map(O => clkfbin3, I => clkfbout3);

  lock300_1 <= flock1 and fdone1;
  lock300_2 <= flock2 and fdone2;
  lock300_3 <= flock3 and fdone3;

  PLL4 : PLL320 port
  map(mclk_in => MCLK40, RESET => RESET, locked => lock320, CLK320 => clk320, CLK40 => TX_CLK);

  PINCAPT_M40_1 : pin_capt port
  map (pin_in => MCLK1, pin_out => MCLK40_IN1, clk600 => clk600_1, clk600_90 => clk600_90_1, clk300 => clk300_1, str => BC_STR1, ptime => BC_BITS1);
  PINCAPT_M40_2 : pin_capt port
  map (pin_in => MCLK2, pin_out => MCLK40_IN2, clk600 => clk600_2, clk600_90 => clk600_90_2, clk300 => clk300_2, str => BC_STR2, ptime => BC_BITS2);
  PINCAPT_M40_3 : pin_capt port
  map (pin_in => MCLK3, pin_out => MCLK40_IN3, clk600 => clk600_3, clk600_90 => clk600_90_3, clk300 => clk300_3, str => BC_STR3, ptime => BC_BITS3);

  TDC1_CHA : TDCCHAN port
  map(pin_in => CGE1i, pin_out => CGE1, clk300 => clk300_1, clk600 => clk600_1, clk600_90 => clk600_90_1, reset => sreset, tdcclk => tdcclk1, rstr => rsa1, rdata => rda1, tdc_count => TDC_COU1, bc_time => BC_PER1, tdc_out => TDC1A, tdc_rdy => TDC1A_rdy0,
  tdc_raw => TDC1A_raw, tdc_raw_lock => spi_lock_1);
  TDC1_CHB : TDCCHAN port
  map(pin_in => CGE2i, pin_out => CGE2, clk300 => clk300_1, clk600 => clk600_1, clk600_90 => clk600_90_1, reset => sreset, tdcclk => tdcclk1, rstr => rsb1, rdata => rdb1, tdc_count => TDC_COU1, bc_time => BC_PER1, tdc_out => TDC1B, tdc_rdy => TDC1B_rdy0,
  tdc_raw => TDC1B_raw, tdc_raw_lock => spi_lock_1);
  TDC1_CHC : TDCCHAN port
  map(pin_in => CGE3i, pin_out => CGE3, clk300 => clk300_1, clk600 => clk600_1, clk600_90 => clk600_90_1, reset => sreset, tdcclk => tdcclk1, rstr => rsc1, rdata => rdc1, tdc_count => TDC_COU1, bc_time => BC_PER1, tdc_out => TDC1C, tdc_rdy => TDC1C_rdy0,
  tdc_raw => TDC1C_raw, tdc_raw_lock => spi_lock_1);
  TDC1_CHD : TDCCHAN port
  map(pin_in => CGE4i, pin_out => CGE4, clk300 => clk300_1, clk600 => clk600_1, clk600_90 => clk600_90_1, reset => sreset, tdcclk => tdcclk1, rstr => rsd1, rdata => rdd1, tdc_count => TDC_COU1, bc_time => BC_PER1, tdc_out => TDC1D, tdc_rdy => TDC1D_rdy0,
  tdc_raw => TDC1D_raw, tdc_raw_lock => spi_lock_1);

  TDC2_CHA : TDCCHAN port
  map(pin_in => CGE5i, pin_out => CGE5, clk300 => clk300_2, clk600 => clk600_2, clk600_90 => clk600_90_2, reset => sreset, tdcclk => tdcclk2, rstr => rsa2, rdata => rda2, tdc_count => TDC_COU2, bc_time => BC_PER2, tdc_out => TDC2A, tdc_rdy => TDC2A_rdy0,
  tdc_raw => TDC2A_raw, tdc_raw_lock => spi_lock_2);
  TDC2_CHB : TDCCHAN port
  map(pin_in => CGE6i, pin_out => CGE6, clk300 => clk300_2, clk600 => clk600_2, clk600_90 => clk600_90_2, reset => sreset, tdcclk => tdcclk2, rstr => rsb2, rdata => rdb2, tdc_count => TDC_COU2, bc_time => BC_PER2, tdc_out => TDC2B, tdc_rdy => TDC2B_rdy0,
  tdc_raw => TDC2B_raw, tdc_raw_lock => spi_lock_2);
  TDC2_CHC : TDCCHAN port
  map(pin_in => CGE7i, pin_out => CGE7, clk300 => clk300_2, clk600 => clk600_2, clk600_90 => clk600_90_2, reset => sreset, tdcclk => tdcclk2, rstr => rsc2, rdata => rdc2, tdc_count => TDC_COU2, bc_time => BC_PER2, tdc_out => TDC2C, tdc_rdy => TDC2C_rdy0,
  tdc_raw => TDC2C_raw, tdc_raw_lock => spi_lock_2);
  TDC2_CHD : TDCCHAN port
  map(pin_in => CGE8i, pin_out => CGE8, clk300 => clk300_2, clk600 => clk600_2, clk600_90 => clk600_90_2, reset => sreset, tdcclk => tdcclk2, rstr => rsd2, rdata => rdd2, tdc_count => TDC_COU2, bc_time => BC_PER2, tdc_out => TDC2D, tdc_rdy => TDC2D_rdy0,
  tdc_raw => TDC2D_raw, tdc_raw_lock => spi_lock_2);

  TDC3_CHA : TDCCHAN port
  map(pin_in => CGE9i, pin_out => CGE9, clk300 => clk300_3, clk600 => clk600_3, clk600_90 => clk600_90_3, reset => sreset, tdcclk => tdcclk3, rstr => rsa3, rdata => rda3, tdc_count => TDC_COU3, bc_time => BC_PER3, tdc_out => TDC3A, tdc_rdy => TDC3A_rdy0,
  tdc_raw => TDC3A_raw, tdc_raw_lock => spi_lock_3);
  TDC3_CHB : TDCCHAN port
  map(pin_in => CGE10i, pin_out => CGE10, clk300 => clk300_3, clk600 => clk600_3, clk600_90 => clk600_90_3, reset => sreset, tdcclk => tdcclk3, rstr => rsb3, rdata => rdb3, tdc_count => TDC_COU3, bc_time => BC_PER3, tdc_out => TDC3B, tdc_rdy => TDC3B_rdy0,
  tdc_raw => TDC3B_raw, tdc_raw_lock => spi_lock_3);
  TDC3_CHC : TDCCHAN port
  map(pin_in => CGE11i, pin_out => CGE11, clk300 => clk300_3, clk600 => clk600_3, clk600_90 => clk600_90_3, reset => sreset, tdcclk => tdcclk3, rstr => rsc3, rdata => rdc3, tdc_count => TDC_COU3, bc_time => BC_PER3, tdc_out => TDC3C, tdc_rdy => TDC3C_rdy0,
  tdc_raw => TDC3C_raw, tdc_raw_lock => spi_lock_3);
  TDC3_CHD : TDCCHAN port
  map(pin_in => CGE12i, pin_out => CGE12, clk300 => clk300_3, clk600 => clk600_3, clk600_90 => clk600_90_3, reset => sreset, tdcclk => tdcclk3, rstr => rsd3, rdata => rdd3, tdc_count => TDC_COU3, bc_time => BC_PER3, tdc_out => TDC3D, tdc_rdy => TDC3D_rdy0,
  tdc_raw => TDC3D_raw, tdc_raw_lock => spi_lock_3);

  CHANNEL1A : channel port
  map (CGE => CGE1, clk320 => clk320, reset => sreset, tdc_rdy_in => TDC1A_rdy0, mt_cou => mt_cou, bc_cou => BC_COU(5 downto 0), TR_bc => TR_to, TDC => TDC1A, CSTR => CSTR1, CH => CH1, CH_shift => CH1A_shift,
  gate_time_low => gate_time_low, gate_time_high => gate_time_high, Ampl_sat => Ampl_sat, ampl_low => ampl_low, CH0_zero => CH1_0_zero, CH1_zero => CH1_1_zero, CH_trig_outt => CH_trig(0), CH_trig_outa => CH_triga(0), CH_trig_bgnd => trig_bgnd(0), CH_TIME => CH_TIME_T(0),
  CH_ampl => CH_ampl0(0), DATA_out => DATA_out(0), DATA_ready => DATA_rdy(0), DATA_rd => DATA_rd(0), FIFO_dis => FIFO_dis, Event_in => Event_in(0), Z0_cal => CH1_Z0, Z1_cal => CH1_Z1, Z_alarm => Z_alarm(0), spi_lock => spi_lock320, R0_cal => CH1_0_rg,
  R1_cal => CH1_1_rg, R0_corr => CH1_0_rc, R1_corr => CH1_1_rc, pulse_in => inp_cou(0), chan_ena => chans_ena(0), trig_dis => trig_dis(0), fdd => fdd, ch_trig_int => ch_trig_outtn(1), ch_trig_outtn => ch_trig_outtn(0));

  CHANNEL1B : channel port
  map (CGE => CGE2, clk320 => clk320, reset => sreset, tdc_rdy_in => TDC1B_rdy0, mt_cou => mt_cou, bc_cou => BC_COU(5 downto 0), TR_bc => TR_to, TDC => TDC1B, CSTR => CSTR2, CH => CH2, CH_shift => CH1B_shift,
  gate_time_low => gate_time_low, gate_time_high => gate_time_high, Ampl_sat => Ampl_sat, ampl_low => ampl_low, CH0_zero => CH2_0_zero, CH1_zero => CH2_1_zero, CH_trig_outt => CH_trig(1), CH_trig_outa => CH_triga(1), CH_trig_bgnd => trig_bgnd(1), CH_TIME => CH_TIME_T(1),
  CH_ampl => CH_ampl0(1), DATA_out => DATA_out(1), DATA_ready => DATA_rdy(1), DATA_rd => DATA_rd(1), FIFO_dis => FIFO_dis, Event_in => Event_in(1), Z0_cal => CH2_Z0, Z1_cal => CH2_Z1, Z_alarm => Z_alarm(1), spi_lock => spi_lock320, R0_cal => CH2_0_rg,
  R1_cal => CH2_1_rg, R0_corr => CH2_0_rc, R1_corr => CH2_1_rc, pulse_in => inp_cou(1), chan_ena => chans_ena(1), trig_dis => trig_dis(1), fdd => fdd, ch_trig_int => ch_trig_outtn(0), ch_trig_outtn => ch_trig_outtn(1));

  CHANNEL1C : channel port
  map (CGE => CGE3, clk320 => clk320, reset => sreset, tdc_rdy_in => TDC1C_rdy0, mt_cou => mt_cou, bc_cou => BC_COU(5 downto 0), TR_bc => TR_to, TDC => TDC1C, CSTR => CSTR3, CH => CH3, CH_shift => CH1C_shift,
  gate_time_low => gate_time_low, gate_time_high => gate_time_high, Ampl_sat => Ampl_sat, ampl_low => ampl_low, CH0_zero => CH3_0_zero, CH1_zero => CH3_1_zero, CH_trig_outt => CH_trig(2), CH_trig_outa => CH_triga(2), CH_trig_bgnd => trig_bgnd(2), CH_TIME => CH_TIME_T(2),
  CH_ampl => CH_ampl0(2), DATA_out => DATA_out(2), DATA_ready => DATA_rdy(2), DATA_rd => DATA_rd(2), FIFO_dis => FIFO_dis, Event_in => Event_in(2), Z0_cal => CH3_Z0, Z1_cal => CH3_Z1, Z_alarm => Z_alarm(2), spi_lock => spi_lock320, R0_cal => CH3_0_rg,
  R1_cal => CH3_1_rg, R0_corr => CH3_0_rc, R1_corr => CH3_1_rc, pulse_in => inp_cou(2), chan_ena => chans_ena(2), trig_dis => trig_dis(2), fdd => fdd, ch_trig_int => ch_trig_outtn(3), ch_trig_outtn => ch_trig_outtn(2));

  CHANNEL1D : channel port
  map (CGE => CGE4, clk320 => clk320, reset => sreset, tdc_rdy_in => TDC1D_rdy0, mt_cou => mt_cou, bc_cou => BC_COU(5 downto 0), TR_bc => TR_to, TDC => TDC1D, CSTR => CSTR4, CH => CH4, CH_shift => CH1D_shift,
  gate_time_low => gate_time_low, gate_time_high => gate_time_high, Ampl_sat => Ampl_sat, ampl_low => ampl_low, CH0_zero => CH4_0_zero, CH1_zero => CH4_1_zero, CH_trig_outt => CH_trig(3), CH_trig_outa => CH_triga(3), CH_trig_bgnd => trig_bgnd(3), CH_TIME => CH_TIME_T(3),
  CH_ampl => CH_ampl0(3), DATA_out => DATA_out(3), DATA_ready => DATA_rdy(3), DATA_rd => DATA_rd(3), FIFO_dis => FIFO_dis, Event_in => Event_in(3), Z0_cal => CH4_Z0, Z1_cal => CH4_Z1, Z_alarm => Z_alarm(3), spi_lock => spi_lock320, R0_cal => CH4_0_rg,
  R1_cal => CH4_1_rg, R0_corr => CH4_0_rc, R1_corr => CH4_1_rc, pulse_in => inp_cou(3), chan_ena => chans_ena(3), trig_dis => trig_dis(3), fdd => fdd, ch_trig_int => ch_trig_outtn(2), ch_trig_outtn => ch_trig_outtn(3));

  CHANNEL2A : channel port
  map (CGE => CGE5, clk320 => clk320, reset => sreset, tdc_rdy_in => TDC2A_rdy0, mt_cou => mt_cou, bc_cou => BC_COU(5 downto 0), TR_bc => TR_to, TDC => TDC2A, CSTR => CSTR5, CH => CH5, CH_shift => CH2A_shift,
  gate_time_low => gate_time_low, gate_time_high => gate_time_high, Ampl_sat => Ampl_sat, ampl_low => ampl_low, CH0_zero => CH5_0_zero, CH1_zero => CH5_1_zero, CH_trig_outt => CH_trig(4), CH_trig_outa => CH_triga(4), CH_trig_bgnd => trig_bgnd(4), CH_TIME => CH_TIME_T(4),
  CH_ampl => CH_ampl0(4), DATA_out => DATA_out(4), DATA_ready => DATA_rdy(4), DATA_rd => DATA_rd(4), FIFO_dis => FIFO_dis, Event_in => Event_in(4), Z0_cal => CH5_Z0, Z1_cal => CH5_Z1, Z_alarm => Z_alarm(4), spi_lock => spi_lock320, R0_cal => CH5_0_rg,
  R1_cal => CH5_1_rg, R0_corr => CH5_0_rc, R1_corr => CH5_1_rc, pulse_in => inp_cou(4), chan_ena => chans_ena(4), trig_dis => trig_dis(4), fdd => fdd, ch_trig_int => ch_trig_outtn(5), ch_trig_outtn => ch_trig_outtn(4));

  CHANNEL2B : channel port
  map (CGE => CGE6, clk320 => clk320, reset => sreset, tdc_rdy_in => TDC2B_rdy0, mt_cou => mt_cou, bc_cou => BC_COU(5 downto 0), TR_bc => TR_to, TDC => TDC2B, CSTR => CSTR6, CH => CH6, CH_shift => CH2B_shift,
  gate_time_low => gate_time_low, gate_time_high => gate_time_high, Ampl_sat => Ampl_sat, ampl_low => ampl_low, CH0_zero => CH6_0_zero, CH1_zero => CH6_1_zero, CH_trig_outt => CH_trig(5), CH_trig_outa => CH_triga(5), CH_trig_bgnd => trig_bgnd(5), CH_TIME => CH_TIME_T(5),
  CH_ampl => CH_ampl0(5), DATA_out => DATA_out(5), DATA_ready => DATA_rdy(5), DATA_rd => DATA_rd(5), FIFO_dis => FIFO_dis, Event_in => Event_in(5), Z0_cal => CH6_Z0, Z1_cal => CH6_Z1, Z_alarm => Z_alarm(5), spi_lock => spi_lock320, R0_cal => CH6_0_rg,
  R1_cal => CH6_1_rg, R0_corr => CH6_0_rc, R1_corr => CH6_1_rc, pulse_in => inp_cou(5), chan_ena => chans_ena(5), trig_dis => trig_dis(5), fdd => fdd, ch_trig_int => ch_trig_outtn(4), ch_trig_outtn => ch_trig_outtn(5));

  CHANNEL2C : channel port
  map (CGE => CGE7, clk320 => clk320, reset => sreset, tdc_rdy_in => TDC2C_rdy0, mt_cou => mt_cou, bc_cou => BC_COU(5 downto 0), TR_bc => TR_to, TDC => TDC2C, CSTR => CSTR7, CH => CH7, CH_shift => CH2C_shift,
  gate_time_low => gate_time_low, gate_time_high => gate_time_high, Ampl_sat => Ampl_sat, ampl_low => ampl_low, CH0_zero => CH7_0_zero, CH1_zero => CH7_1_zero, CH_trig_outt => CH_trig(6), CH_trig_outa => CH_triga(6), CH_trig_bgnd => trig_bgnd(6), CH_TIME => CH_TIME_T(6),
  CH_ampl => CH_ampl0(6), DATA_out => DATA_out(6), DATA_ready => DATA_rdy(6), DATA_rd => DATA_rd(6), FIFO_dis => FIFO_dis, Event_in => Event_in(6), Z0_cal => CH7_Z0, Z1_cal => CH7_Z1, Z_alarm => Z_alarm(6), spi_lock => spi_lock320, R0_cal => CH7_0_rg,
  R1_cal => CH7_1_rg, R0_corr => CH7_0_rc, R1_corr => CH7_1_rc, pulse_in => inp_cou(6), chan_ena => chans_ena(6), trig_dis => trig_dis(6), fdd => fdd, ch_trig_int => ch_trig_outtn(7), ch_trig_outtn => ch_trig_outtn(6));

  CHANNEL2D : channel port
  map (CGE => CGE8, clk320 => clk320, reset => sreset, tdc_rdy_in => TDC2D_rdy0, mt_cou => mt_cou, bc_cou => BC_COU(5 downto 0), TR_bc => TR_to, TDC => TDC2D, CSTR => CSTR8, CH => CH8, CH_shift => CH2D_shift,
  gate_time_low => gate_time_low, gate_time_high => gate_time_high, Ampl_sat => Ampl_sat, ampl_low => ampl_low, CH0_zero => CH8_0_zero, CH1_zero => CH8_1_zero, CH_trig_outt => CH_trig(7), CH_trig_outa => CH_triga(7), CH_trig_bgnd => trig_bgnd(7), CH_TIME => CH_TIME_T(7),
  CH_ampl => CH_ampl0(7), DATA_out => DATA_out(7), DATA_ready => DATA_rdy(7), DATA_rd => DATA_rd(7), FIFO_dis => FIFO_dis, Event_in => Event_in(7), Z0_cal => CH8_Z0, Z1_cal => CH8_Z1, Z_alarm => Z_alarm(7), spi_lock => spi_lock320, R0_cal => CH8_0_rg,
  R1_cal => CH8_1_rg, R0_corr => CH8_0_rc, R1_corr => CH8_1_rc, pulse_in => inp_cou(7), chan_ena => chans_ena(7), trig_dis => trig_dis(7), fdd => fdd, ch_trig_int => ch_trig_outtn(6), ch_trig_outtn => ch_trig_outtn(7));

  CHANNEL3A : channel port
  map (CGE => CGE9, clk320 => clk320, reset => sreset, tdc_rdy_in => TDC3A_rdy0, mt_cou => mt_cou, bc_cou => BC_COU(5 downto 0), TR_bc => TR_to, TDC => TDC3A, CSTR => CSTR9, CH => CH9, CH_shift => CH3A_shift,
  gate_time_low => gate_time_low, gate_time_high => gate_time_high, Ampl_sat => Ampl_sat, ampl_low => ampl_low, CH0_zero => CH9_0_zero, CH1_zero => CH9_1_zero, CH_trig_outt => CH_trig(8), CH_trig_outa => CH_triga(8), CH_trig_bgnd => trig_bgnd(8), CH_TIME => CH_TIME_T(8),
  CH_ampl => CH_ampl0(8), DATA_out => DATA_out(8), DATA_ready => DATA_rdy(8), DATA_rd => DATA_rd(8), FIFO_dis => FIFO_dis, Event_in => Event_in(8), Z0_cal => CH9_Z0, Z1_cal => CH9_Z1, Z_alarm => Z_alarm(8), spi_lock => spi_lock320, R0_cal => CH9_0_rg,
  R1_cal => CH9_1_rg, R0_corr => CH9_0_rc, R1_corr => CH9_1_rc, pulse_in => inp_cou(8), chan_ena => chans_ena(8), trig_dis => trig_dis(8), fdd => fdd, ch_trig_int => ch_trig_outtn(9), ch_trig_outtn => ch_trig_outtn(8));

  CHANNEL3B : channel port
  map (CGE => CGE10, clk320 => clk320, reset => sreset, tdc_rdy_in => TDC3B_rdy0, mt_cou => mt_cou, bc_cou => BC_COU(5 downto 0), TR_bc => TR_to, TDC => TDC3B, CSTR => CSTR10, CH => CH10, CH_shift => CH3B_shift,
  gate_time_low => gate_time_low, gate_time_high => gate_time_high, Ampl_sat => Ampl_sat, ampl_low => ampl_low, CH0_zero => CH10_0_zero, CH1_zero => CH10_1_zero, CH_trig_outt => CH_trig(9), CH_trig_outa => CH_triga(9), CH_trig_bgnd => trig_bgnd(9), CH_TIME => CH_TIME_T(9),
  CH_ampl => CH_ampl0(9), DATA_out => DATA_out(9), DATA_ready => DATA_rdy(9), DATA_rd => DATA_rd(9), FIFO_dis => FIFO_dis, Event_in => Event_in(9), Z0_cal => CH10_Z0, Z1_cal => CH10_Z1, Z_alarm => Z_alarm(9), spi_lock => spi_lock320, R0_cal => CH10_0_rg,
  R1_cal => CH10_1_rg, R0_corr => CH10_0_rc, R1_corr => CH10_1_rc, pulse_in => inp_cou(9), chan_ena => chans_ena(9), trig_dis => trig_dis(9), fdd => fdd, ch_trig_int => ch_trig_outtn(8), ch_trig_outtn => ch_trig_outtn(9));

  CHANNEL3C : channel port
  map (CGE => CGE11, clk320 => clk320, reset => sreset, tdc_rdy_in => TDC3C_rdy0, mt_cou => mt_cou, bc_cou => BC_COU(5 downto 0), TR_bc => TR_to, TDC => TDC3C, CSTR => CSTR11, CH => CH11, CH_shift => CH3C_shift,
  gate_time_low => gate_time_low, gate_time_high => gate_time_high, Ampl_sat => Ampl_sat, ampl_low => ampl_low, CH0_zero => CH11_0_zero, CH1_zero => CH11_1_zero, CH_trig_outt => CH_trig(10), CH_trig_outa => CH_triga(10), CH_trig_bgnd => trig_bgnd(10), CH_TIME => CH_TIME_T(10),
  CH_ampl => CH_ampl0(10), DATA_out => DATA_out(10), DATA_ready => DATA_rdy(10), DATA_rd => DATA_rd(10), FIFO_dis => FIFO_dis, Event_in => Event_in(10), Z0_cal => CH11_Z0, Z1_cal => CH11_Z1, Z_alarm => Z_alarm(10), spi_lock => spi_lock320, R0_cal => CH11_0_rg,
  R1_cal => CH11_1_rg, R0_corr => CH11_0_rc, R1_corr => CH11_1_rc, pulse_in => inp_cou(10), chan_ena => chans_ena(10), trig_dis => trig_dis(10), fdd => fdd, ch_trig_int => ch_trig_outtn(11), ch_trig_outtn => ch_trig_outtn(10));

  CHANNEL3D : channel port
  map (CGE => CGE12, clk320 => clk320, reset => sreset, tdc_rdy_in => TDC3D_rdy0, mt_cou => mt_cou, bc_cou => BC_COU(5 downto 0), TR_bc => TR_to, TDC => TDC3D, CSTR => CSTR12, CH => CH12, CH_shift => CH3D_shift,
  gate_time_low => gate_time_low, gate_time_high => gate_time_high, Ampl_sat => Ampl_sat, ampl_low => ampl_low, CH0_zero => CH12_0_zero, CH1_zero => CH12_1_zero, CH_trig_outt => CH_trig(11), CH_trig_outa => CH_triga(11), CH_trig_bgnd => trig_bgnd(11), CH_TIME => CH_TIME_T(11),
  CH_ampl => CH_ampl0(11), DATA_out => DATA_out(11), DATA_ready => DATA_rdy(11), DATA_rd => DATA_rd(11), FIFO_dis => FIFO_dis, Event_in => Event_in(11), Z0_cal => CH12_Z0, Z1_cal => CH12_Z1, Z_alarm => Z_alarm(11), spi_lock => spi_lock320, R0_cal => CH12_0_rg,
  R1_cal => CH12_1_rg, R0_corr => CH12_0_rc, R1_corr => CH12_1_rc, pulse_in => inp_cou(11), chan_ena => chans_ena(11), trig_dis => trig_dis(11), fdd => fdd, ch_trig_int => ch_trig_outtn(10), ch_trig_outtn => ch_trig_outtn(11));

  TRG0 : trigger port
  map (clk320 => clk320, mt_cou => mt_cou, CH_trigt => CH_trig, CH_triga => CH_triga, CH_trigb => trig_bgnd, CH_TIME_T => CH_TIME_T, CH_ampl0 => CH_ampl0, tcm_req => tcm_req, tt => tt, ta => ta);

  EV_FIFO : EVENTID_FIFO port
  map (clk => clk320, srst => sreset, din => EV_ID_in, wr_en => EV_ID_wr, rd_en => EV_ID_rd, dout => EV_ID_out, full => open, empty => EV_ID_empty);

  EV_ID_in <= Orbit_ID & BC_Cou & Event_in;
  EV_ID_wr <= '1' when (inp_event = '1') and (mt_cou = "001") else
    '0';
  EV_ID_rd <= '1' when (EV_ID_empty = '0') and ((Event_free = '1') or ((Event_ready = '1') and (CH_do = 0)) or (ev_tout = '1')) else
    '0';

  --OUT_FIFO: FIFO_OUT port map (rst =>sreset, wr_clk => clk320, rd_clk=>TX_CLK, din =>DATA80_in, wr_en => WR_fifo_out, rd_en =>DATA80_rd, dout => DATA80_out, full =>open, empty =>DATA_empty, wr_rst_busy => open, rd_rst_busy => open);

  --DATA80_rd<= not DATA_empty;

  count1 : counters port
  map (clk => clk320, evnt => inp_cou, trig => cnt_trig, reset => cnt_rst, dout => cnt_out, hdout => hcnt_out, raddr => spi_addr(5 downto 0), hraddr => hspi_addr(4 downto 0), hl => hspi_h, rd_en => cnt_rd, hrd_en => hcnt_rd);

  process (MCLK40, RESET)
  begin
    if (RESET = '1') then
      sreset   <= '1';
      rstcount <= "0000";
    else
      if (MCLK40'event) and (MCLK40 = '1') then

        alm_rst0   <= sreset;
        all_locked <= lock320 and lock300_1 and lock300_2 and lock300_3;

        if (rstcount = "1111") then
          sreset <= '0';
        else
          if (all_locked = '1') then
            rstcount <= rstcount + 1;
          end if;
        end if;
      end if;
    end if;
  end process;

  alm_rst <= not sreset and alm_rst0;

  rd_lock_hspi <= '1' when (hspi_bit_count(3 downto 0) = x"F") and (hspi_rd = '1') and (hspi_addr(8) = '0') else
    '0';
  Hs_rd <= alm_rst or Hs_clr;

  flsh_sel <= '1' when (hspi_addr(7 downto 2) = "111110") else
    '0';
  rdo_sel <= '1' when (hspi_addr >= 16#E8#) and (hspi_addr <= 16#F4#) else
    '0';
  rd_xadc <= '1' when (hspi_addr >= 16#FC#) and (hspi_addr <= 16#FE#) else
    '0';
  hysta_sel <= '1' when (hspi_addr = 16#F5#) else
    '0';
  hystd_sel <= '1' when (hspi_addr = 16#F6#) else
    '0';

  process (HSCKI, HSELI, RESET)
  begin
    if (HSELI = '0') then
      hspi_bit_count <= "00000";
      hcnt_rd        <= '0';
      hspibuf_wr     <= '0';
      hspibuf_rd     <= '0';
      hspi_na        <= '0';
      reg32_wr       <= '0';
      Hs_clr         <= '0';
      reg32_rd       <= '0';
      reg32_str      <= '0';
    else

      if (HSCKI'event and HSCKI = '0') then

        if (hspi_bit_count = "11111") then
          hspi_bit_count <= "10000";
          hspi_na        <= '1';
          if (hspi_rd = '0') then
            if (hspi_h = '0') then
              hspi_wr_data <= HSPI_DATA(14 downto 0) & HMOSII;
            else
              hspi_wr_data_l <= HSPI_DATA(14 downto 0) & HMOSII;
            end if;
            if (hspi_addr(7) = '0') then
              hspi_wr_rdy <= '1';
            end if;
            if (hspi_addr(7 downto 6) = "10") and (hspi_addr(5 downto 2) /= "1111") then
              hspibuf_wr <= '1';
            end if;
            if (hspi_addr(7 downto 3) >= "11011") and (hspi_h = '1') then
              reg32_wr <= '1';
            end if;

          end if;
        else
          hspi_bit_count <= hspi_bit_count + 1;
        end if;

        if (hspi_bit_count = "10000") then
          hspi_wr_rdy <= '0';
          hspibuf_wr  <= '0';
          reg32_wr    <= '0';
          if (hspi_rd = '0') and (hspi_na = '1') then
            if (hspi_addr(7 downto 4) < x"C") or (hspi_h = '1') then
              hspi_addr <= hspi_addr + 1;
            end if;
            if (hspi_addr(7 downto 3) >= "11011") then
              hspi_h <= not hspi_h;
            end if;
          end if;
        end if;

        if ((hspi_bit_count = "01010") or ((hspi_bit_count = "10001") and (hspi_h = '0'))) and (hspi_rd = '1') then
          reg32_rd <= '1';
        else
          reg32_rd <= '0';
        end if;

        if (hspi_bit_count = "10001") and (hspi_h = '1') and (hspi_rd = '1') then
          reg32_str <= '1';
        else
          reg32_str <= '0';
        end if;
        if (hspi_bit_count = "10001") and (hspi_rd = '1') and (hspi_addr = 16#80#) then
          Hs_clr <= '1';
        else
          Hs_clr <= '0';
        end if;

        if (hspi_bit_count = "00000") then
          hspi_rd <= HMOSII;
        end if;
        if (hspi_bit_count = "01001") then
          hspi_addr <= HSPI_DATA(7 downto 0) & HMOSII;
          hspi_h    <= '0';
        end if;
        if (hspi_bit_count = "01110") and (hspi_rd = '1') and (hspi_addr(7 downto 0) = x"C0") then
          hcnt_rd <= '1';
        end if;

        if (hspi_bit_count(3 downto 0) = "1110") and (hspi_rd = '1') and (hspi_addr(7 downto 6) = "10") then
          hspibuf_rd <= '1';
        end if;

        if (rd_lock_hspi = '1') then
          hspibuf_rd <= '0';

          if (hspi_addr(7 downto 4) >= x"C") then
            hspi_h <= not hspi_h;
          end if;
          if ((hspi_addr(7 downto 4) < x"C") or (hspi_h = '1')) then
            hspi_addr <= hspi_addr + 1;
          end if;
          if (hspi_addr(7 downto 3) >= "11011") and (hspi_h = '1') then
            HSPI_DATA <= hspi_32l;

          else

            case to_integer(unsigned(hspi_addr(7 downto 0))) is
              when 0     => HSPI_DATA     <= "0000000" & fdd & gate_time_high;
              when 1     => HSPI_DATA     <= "000" & trig_dis(0) & CH1A_shift;
              when 2     => HSPI_DATA     <= "000" & trig_dis(1) & CH1B_shift;
              when 3     => HSPI_DATA     <= "000" & trig_dis(2) & CH1C_shift;
              when 4     => HSPI_DATA     <= "000" & trig_dis(3) & CH1D_shift;
              when 5     => HSPI_DATA     <= "000" & trig_dis(4) & CH2A_shift;
              when 6     => HSPI_DATA     <= "000" & trig_dis(5) & CH2B_shift;
              when 7     => HSPI_DATA     <= "000" & trig_dis(6) & CH2C_shift;
              when 8     => HSPI_DATA     <= "000" & trig_dis(7) & CH2D_shift;
              when 9     => HSPI_DATA     <= "000" & trig_dis(8) & CH3A_shift;
              when 16#A# => HSPI_DATA <= "000" & trig_dis(9) & CH3B_shift;
              when 16#B# => HSPI_DATA <= "000" & trig_dis(10) & CH3C_shift;
              when 16#C# => HSPI_DATA <= "000" & trig_dis(11) & CH3D_shift;

              when 16#D#  => HSPI_DATA  <= x"0" & CH1_0_zero;
              when 16#E#  => HSPI_DATA  <= x"0" & CH1_1_zero;
              when 16#F#  => HSPI_DATA  <= x"0" & CH2_0_zero;
              when 16#10# => HSPI_DATA <= x"0" & CH2_1_zero;
              when 16#11# => HSPI_DATA <= x"0" & CH3_0_zero;
              when 16#12# => HSPI_DATA <= x"0" & CH3_1_zero;
              when 16#13# => HSPI_DATA <= x"0" & CH4_0_zero;
              when 16#14# => HSPI_DATA <= x"0" & CH4_1_zero;
              when 16#15# => HSPI_DATA <= x"0" & CH5_0_zero;
              when 16#16# => HSPI_DATA <= x"0" & CH5_1_zero;
              when 16#17# => HSPI_DATA <= x"0" & CH6_0_zero;
              when 16#18# => HSPI_DATA <= x"0" & CH6_1_zero;
              when 16#19# => HSPI_DATA <= x"0" & CH7_0_zero;
              when 16#1A# => HSPI_DATA <= x"0" & CH7_1_zero;
              when 16#1B# => HSPI_DATA <= x"0" & CH8_0_zero;
              when 16#1C# => HSPI_DATA <= x"0" & CH8_1_zero;
              when 16#1D# => HSPI_DATA <= x"0" & CH9_0_zero;
              when 16#1E# => HSPI_DATA <= x"0" & CH9_1_zero;
              when 16#1F# => HSPI_DATA <= x"0" & CH10_0_zero;
              when 16#20# => HSPI_DATA <= x"0" & CH10_1_zero;
              when 16#21# => HSPI_DATA <= x"0" & CH11_0_zero;
              when 16#22# => HSPI_DATA <= x"0" & CH11_1_zero;
              when 16#23# => HSPI_DATA <= x"0" & CH12_0_zero;
              when 16#24# => HSPI_DATA <= x"0" & CH12_1_zero;

              when 16#25# => HSPI_DATA <= x"0" & CH1_0_rc;
              when 16#26# => HSPI_DATA <= x"0" & CH1_1_rc;
              when 16#27# => HSPI_DATA <= x"0" & CH2_0_rc;
              when 16#28# => HSPI_DATA <= x"0" & CH2_1_rc;
              when 16#29# => HSPI_DATA <= x"0" & CH3_0_rc;
              when 16#2A# => HSPI_DATA <= x"0" & CH3_1_rc;
              when 16#2B# => HSPI_DATA <= x"0" & CH4_0_rc;
              when 16#2C# => HSPI_DATA <= x"0" & CH4_1_rc;
              when 16#2D# => HSPI_DATA <= x"0" & CH5_0_rc;
              when 16#2E# => HSPI_DATA <= x"0" & CH5_1_rc;
              when 16#2F# => HSPI_DATA <= x"0" & CH6_0_rc;
              when 16#30# => HSPI_DATA <= x"0" & CH6_1_rc;
              when 16#31# => HSPI_DATA <= x"0" & CH7_0_rc;
              when 16#32# => HSPI_DATA <= x"0" & CH7_1_rc;
              when 16#33# => HSPI_DATA <= x"0" & CH8_0_rc;
              when 16#34# => HSPI_DATA <= x"0" & CH8_1_rc;
              when 16#35# => HSPI_DATA <= x"0" & CH9_0_rc;
              when 16#36# => HSPI_DATA <= x"0" & CH9_1_rc;
              when 16#37# => HSPI_DATA <= x"0" & CH10_0_rc;
              when 16#38# => HSPI_DATA <= x"0" & CH10_1_rc;
              when 16#39# => HSPI_DATA <= x"0" & CH11_0_rc;
              when 16#3A# => HSPI_DATA <= x"0" & CH11_1_rc;
              when 16#3B# => HSPI_DATA <= x"0" & CH12_0_rc;
              when 16#3C# => HSPI_DATA <= x"0" & CH12_1_rc;
              when 16#3D# => HSPI_DATA <= ampl_low & Ampl_sat;

              when 16#3E# => HSPI_DATA <= pshift2(5) & pshift2(5) & pshift2 & pshift1(5) & pshift1(5) & pshift1;
              when 16#3F# => HSPI_DATA <= x"00" & pshift3(5) & pshift3(5) & pshift3;
              when 16#40# => HSPI_DATA <= "00" & TDC1A_raw (12 downto 7) & '0' & TDC1A_raw(6 downto 0);
              when 16#41# => HSPI_DATA <= "00" & TDC1B_raw (12 downto 7) & '0' & TDC1B_raw(6 downto 0);
              when 16#42# => HSPI_DATA <= "00" & TDC1C_raw (12 downto 7) & '0' & TDC1C_raw(6 downto 0);
              when 16#43# => HSPI_DATA <= "00" & TDC1D_raw (12 downto 7) & '0' & TDC1D_raw(6 downto 0);
              when 16#44# => HSPI_DATA <= "00" & TDC2A_raw (12 downto 7) & '0' & TDC2A_raw(6 downto 0);
              when 16#45# => HSPI_DATA <= "00" & TDC2B_raw (12 downto 7) & '0' & TDC2B_raw(6 downto 0);
              when 16#46# => HSPI_DATA <= "00" & TDC2C_raw (12 downto 7) & '0' & TDC2C_raw(6 downto 0);
              when 16#47# => HSPI_DATA <= "00" & TDC2D_raw (12 downto 7) & '0' & TDC2D_raw(6 downto 0);
              when 16#48# => HSPI_DATA <= "00" & TDC3A_raw (12 downto 7) & '0' & TDC3A_raw(6 downto 0);
              when 16#49# => HSPI_DATA <= "00" & TDC3B_raw (12 downto 7) & '0' & TDC3B_raw(6 downto 0);
              when 16#4A# => HSPI_DATA <= "00" & TDC3C_raw (12 downto 7) & '0' & TDC3C_raw(6 downto 0);
              when 16#4B# => HSPI_DATA <= "00" & TDC3D_raw (12 downto 7) & '0' & TDC3D_raw(6 downto 0);

              when 16#4C# => HSPI_DATA <= CH1_Z0;
              when 16#4D# => HSPI_DATA <= CH1_Z1;
              when 16#4E# => HSPI_DATA <= CH2_Z0;
              when 16#4F# => HSPI_DATA <= CH2_Z1;
              when 16#50# => HSPI_DATA <= CH3_Z0;
              when 16#51# => HSPI_DATA <= CH3_Z1;
              when 16#52# => HSPI_DATA <= CH4_Z0;
              when 16#53# => HSPI_DATA <= CH4_Z1;
              when 16#54# => HSPI_DATA <= CH5_Z0;
              when 16#55# => HSPI_DATA <= CH5_Z1;
              when 16#56# => HSPI_DATA <= CH6_Z0;
              when 16#57# => HSPI_DATA <= CH6_Z1;
              when 16#58# => HSPI_DATA <= CH7_Z0;
              when 16#59# => HSPI_DATA <= CH7_Z1;
              when 16#5A# => HSPI_DATA <= CH8_Z0;
              when 16#5B# => HSPI_DATA <= CH8_Z1;
              when 16#5C# => HSPI_DATA <= CH9_Z0;
              when 16#5D# => HSPI_DATA <= CH9_Z1;
              when 16#5E# => HSPI_DATA <= CH10_Z0;
              when 16#5F# => HSPI_DATA <= CH10_Z1;
              when 16#60# => HSPI_DATA <= CH11_Z0;
              when 16#61# => HSPI_DATA <= CH11_Z1;
              when 16#62# => HSPI_DATA <= CH12_Z0;
              when 16#63# => HSPI_DATA <= CH12_Z1;

              when 16#64# => HSPI_DATA <= std_logic_vector(resize(signed(CH1_0_rg), 16));
              when 16#65# => HSPI_DATA <= std_logic_vector(resize(signed(CH1_1_rg), 16));
              when 16#66# => HSPI_DATA <= std_logic_vector(resize(signed(CH2_0_rg), 16));
              when 16#67# => HSPI_DATA <= std_logic_vector(resize(signed(CH2_1_rg), 16));
              when 16#68# => HSPI_DATA <= std_logic_vector(resize(signed(CH3_0_rg), 16));
              when 16#69# => HSPI_DATA <= std_logic_vector(resize(signed(CH3_1_rg), 16));
              when 16#6A# => HSPI_DATA <= std_logic_vector(resize(signed(CH4_0_rg), 16));
              when 16#6B# => HSPI_DATA <= std_logic_vector(resize(signed(CH4_1_rg), 16));
              when 16#6C# => HSPI_DATA <= std_logic_vector(resize(signed(CH5_0_rg), 16));
              when 16#6D# => HSPI_DATA <= std_logic_vector(resize(signed(CH5_1_rg), 16));
              when 16#6E# => HSPI_DATA <= std_logic_vector(resize(signed(CH6_0_rg), 16));
              when 16#6F# => HSPI_DATA <= std_logic_vector(resize(signed(CH6_1_rg), 16));
              when 16#70# => HSPI_DATA <= std_logic_vector(resize(signed(CH7_0_rg), 16));
              when 16#71# => HSPI_DATA <= std_logic_vector(resize(signed(CH7_1_rg), 16));
              when 16#72# => HSPI_DATA <= std_logic_vector(resize(signed(CH8_0_rg), 16));
              when 16#73# => HSPI_DATA <= std_logic_vector(resize(signed(CH8_1_rg), 16));
              when 16#74# => HSPI_DATA <= std_logic_vector(resize(signed(CH9_0_rg), 16));
              when 16#75# => HSPI_DATA <= std_logic_vector(resize(signed(CH9_1_rg), 16));
              when 16#76# => HSPI_DATA <= std_logic_vector(resize(signed(CH10_0_rg), 16));
              when 16#77# => HSPI_DATA <= std_logic_vector(resize(signed(CH10_1_rg), 16));
              when 16#78# => HSPI_DATA <= std_logic_vector(resize(signed(CH11_0_rg), 16));
              when 16#79# => HSPI_DATA <= std_logic_vector(resize(signed(CH11_1_rg), 16));
              when 16#7A# => HSPI_DATA <= std_logic_vector(resize(signed(CH12_0_rg), 16));
              when 16#7B# => HSPI_DATA <= std_logic_vector(resize(signed(CH12_1_rg), 16));

              when 16#7C#           => HSPI_DATA           <= x"0" & chans_ena_r;
              when 16#7D#           => HSPI_DATA           <= x"0" & Z_alarm;
              when 16#7E#           => HSPI_DATA           <= hyst_md;
              when 16#7F#           => HSPI_DATA           <= gbt_global_status & is_rst & cnt_md & h_busy & HBC_JUMP3 & HBC_JUMP2 & HBC_JUMP1 & HGBTRXerr & GBTRX_ready & lock300_3 & lock300_2 & lock300_1 & lock320;
              when 16#80# to 16#BF# => HSPI_DATA <= hspi_buf_out;

              when 16#C0# to 16#D7# => HSPI_DATA <= hcnt_out;

                -- gbt status            ipbus_control_reg
              when 16#D8# to 16#e7# => HSPI_DATA <= ipbus_control_reg(to_integer(unsigned(hspi_addr(7 downto 0))) - 16#D8#)(31 downto 16);
                hspi_32l                           <= ipbus_control_reg(to_integer(unsigned(hspi_addr(7 downto 0))) - 16#D8#)(15 downto 0);

              when 16#E8# to 16#F4# =>
                HSPI_DATA <= hspib_32(31 downto 16);
                hspi_32l  <= hspib_32(15 downto 0);

              when 16#F5# =>
                HSPI_DATA <= x"000" & "000" & hyst_addr(16);
                hspi_32l  <= hyst_addr(15 downto 0);

              when 16#F6# =>
                HSPI_DATA <= hyst_r_data(31 downto 16);
                hspi_32l  <= hyst_r_data(15 downto 0);

              when 16#F7# => HSPI_DATA <= mcu_tstamp(31 downto 16);
                hspi_32l                 <= mcu_tstamp(15 downto 0);

              when 16#F8# to 16#FB# => HSPI_DATA <= hspib_32(31 downto 16);
                hspi_32l                           <= hspib_32(15 downto 0);

              when 16#FC# to 16#FE# => HSPI_DATA <= (others => '0');
                hspi_32l                           <= xadc_r;

              when 16#FF# => HSPI_DATA <= tstamp(31 downto 16);
                hspi_32l                 <= tstamp(15 downto 0);
              when others => HSPI_DATA <= x"0000";

            end case;
          end if;
        else
          HSPI_DATA <= HSPI_DATA(14 downto 0) & HMOSII;
        end if;

      end if;
    end if;
  end process;

  h0 : hyst port
  map(clk320 => clk320, hyst_inp_data => hyst_data, hyst_a => hyst_a, hyst_t => hyst_t, hyst_st => start_hyst, cnt_clr => hyst_clr, busy => h_busy, hyst_addr_i => hspid_w32(16 downto 0), hyst_addr_o => hyst_addr,
  wr_addr => wr_hyst_a, hyst_data_o => hyst_r_data, n_addr => rd_hyst_d, lock320 => hspi_lock320, stp => hyst_stp);

  wr_hyst_a <= reg32_320_wr and hysta_sel;
  rd_hyst_d <= reg32_320_str and hystd_sel;
  hyst_clr  <= cnt_rst or hyst_rst;

  h1 : for i in 0 to 11 generate
    hyst_data(i) <= DATA_out(i)(25 downto 0);
    hyst_a(i)    <= EV_ID_out(i) and DATA_out(i)(28);
    hyst_t(i)    <= EV_ID_out(i) and not (DATA_out(i)(27) or DATA_out(i)(32));
  end generate;
  UA2 : USR_ACCESSE2 port
  map (CFGCLK => open, DATA => tstamp, DATAVALID => open);

  SNS : SENSOR port
  map (di_in => (others => '0'), daddr_in => xadc_a, den_in => xadc_en, dwe_in => '0', drdy_out => xadc_rdy, do_out => xadc_out, dclk_in => TX_CLK,
  reset_in => sreset, vp_in => '0', vn_in => '0', channel_out => open, eoc_out => open, alarm_out => open, eos_out => open, busy_out => open);

  xadc_a  <= "00000" & hspi_addr(1 downto 0);
  xadc_en <= rd_hspi32 and rd_xadc;

  TCM_reqh <= HBC_JUMP3 or HBC_JUMP2 or HBC_JUMP1 or HGBTRXerr or HGBT_chg;

  rd_lock_spi <= '1' when (spi_bit_count(3 downto 0) = x"F") and (spi_rd = '1') and (spi_addr(8) = '0') else
    '0';
  ALM_CLR <= '1' when (spi_bit_count = "10000") and (spi_rd = '1') and (spi_addr = '0' & x"80") else
    '0';
  buf_lock <= '1' when (spi_bit_count(3 downto 0) = x"A") and (spi_rd = '1') and (spi_addr = '0' & x"F0") else
    '0';

  process (SCKI, SPI_CS)
  begin
    if (SPI_CS = '1') then
      spi_bit_count <= "00000";
      cnt_rd        <= '0';
      spibuf_wr     <= '0';
      spibuf_rd     <= '0';
      spi_na        <= '0';
    else
      if (SCKi'event and SCKi = '0') then
        MISOI <= SPI_DATA(15);
      end if;

      if (SCKI'event and SCKI = '1') then
        if (spi_bit_count = "11111") then
          spi_bit_count <= "10000";
          spi_na        <= '1';
          if (spi_rd = '0') then
            if (spi_addr(7 downto 0) = x"F5") then
              mcu_tstamp(15 downto 0) <= SPI_DATA(14 downto 0) & MOSII;
            end if;
            if (spi_addr(7 downto 0) = x"F6") then
              mcu_tstamp(31 downto 16) <= SPI_DATA(14 downto 0) & MOSII;
            end if;
            spi_wr_data <= SPI_DATA(14 downto 0) & MOSII;
            if (spi_addr(7) = '0') then
              spi_wr_rdy <= '1';
            else
              if (spi_addr(6) = '0') then
                spibuf_wr <= '1';
              end if;
            end if;
          end if;
        else
          spi_bit_count <= spi_bit_count + 1;
        end if;

        if (spi_bit_count = "10000") then
          spi_wr_rdy <= '0';
          spibuf_wr  <= '0';
          if (spi_rd = '0') and (spi_na = '1') then
            spi_addr <= spi_addr + 1;
          end if;
        end if;
        if (spi_bit_count = "00000") then
          spi_rd <= MOSII;
        end if;
        if (spi_bit_count = "01001") then
          spi_addr <= SPI_DATA(7 downto 0) & MOSII;
        end if;
        if (spi_bit_count = "01110") and (spi_rd = '1') and (spi_addr(7 downto 0) = x"C0") then
          cnt_rd <= '1';
        end if;

        if (spi_bit_count(3 downto 0) = "1110") and (spi_rd = '1') and (spi_addr(7 downto 6) = "10") then
          spibuf_rd <= '1';
        end if;

        if (rd_lock_spi = '1') then
          spibuf_rd <= '0';
          spi_addr  <= spi_addr + 1;

          case to_integer(unsigned(spi_addr(7 downto 0))) is
            when 0     => SPI_DATA     <= x"00" & gate_time_high;
            when 1     => SPI_DATA     <= x"0" & CH1A_shift;
            when 2     => SPI_DATA     <= x"0" & CH1B_shift;
            when 3     => SPI_DATA     <= x"0" & CH1C_shift;
            when 4     => SPI_DATA     <= x"0" & CH1D_shift;
            when 5     => SPI_DATA     <= x"0" & CH2A_shift;
            when 6     => SPI_DATA     <= x"0" & CH2B_shift;
            when 7     => SPI_DATA     <= x"0" & CH2C_shift;
            when 8     => SPI_DATA     <= x"0" & CH2D_shift;
            when 9     => SPI_DATA     <= x"0" & CH3A_shift;
            when 16#A# => SPI_DATA <= x"0" & CH3B_shift;
            when 16#B# => SPI_DATA <= x"0" & CH3C_shift;
            when 16#C# => SPI_DATA <= x"0" & CH3D_shift;

            when 16#D#  => SPI_DATA  <= x"0" & CH1_0_zero;
            when 16#E#  => SPI_DATA  <= x"0" & CH1_1_zero;
            when 16#F#  => SPI_DATA  <= x"0" & CH2_0_zero;
            when 16#10# => SPI_DATA <= x"0" & CH2_1_zero;
            when 16#11# => SPI_DATA <= x"0" & CH3_0_zero;
            when 16#12# => SPI_DATA <= x"0" & CH3_1_zero;
            when 16#13# => SPI_DATA <= x"0" & CH4_0_zero;
            when 16#14# => SPI_DATA <= x"0" & CH4_1_zero;
            when 16#15# => SPI_DATA <= x"0" & CH5_0_zero;
            when 16#16# => SPI_DATA <= x"0" & CH5_1_zero;
            when 16#17# => SPI_DATA <= x"0" & CH6_0_zero;
            when 16#18# => SPI_DATA <= x"0" & CH6_1_zero;
            when 16#19# => SPI_DATA <= x"0" & CH7_0_zero;
            when 16#1A# => SPI_DATA <= x"0" & CH7_1_zero;
            when 16#1B# => SPI_DATA <= x"0" & CH8_0_zero;
            when 16#1C# => SPI_DATA <= x"0" & CH8_1_zero;
            when 16#1D# => SPI_DATA <= x"0" & CH9_0_zero;
            when 16#1E# => SPI_DATA <= x"0" & CH9_1_zero;
            when 16#1F# => SPI_DATA <= x"0" & CH10_0_zero;
            when 16#20# => SPI_DATA <= x"0" & CH10_1_zero;
            when 16#21# => SPI_DATA <= x"0" & CH11_0_zero;
            when 16#22# => SPI_DATA <= x"0" & CH11_1_zero;
            when 16#23# => SPI_DATA <= x"0" & CH12_0_zero;
            when 16#24# => SPI_DATA <= x"0" & CH12_1_zero;

            when 16#25# => SPI_DATA <= x"0" & CH1_0_rc;
            when 16#26# => SPI_DATA <= x"0" & CH1_1_rc;
            when 16#27# => SPI_DATA <= x"0" & CH2_0_rc;
            when 16#28# => SPI_DATA <= x"0" & CH2_1_rc;
            when 16#29# => SPI_DATA <= x"0" & CH3_0_rc;
            when 16#2A# => SPI_DATA <= x"0" & CH3_1_rc;
            when 16#2B# => SPI_DATA <= x"0" & CH4_0_rc;
            when 16#2C# => SPI_DATA <= x"0" & CH4_1_rc;
            when 16#2D# => SPI_DATA <= x"0" & CH5_0_rc;
            when 16#2E# => SPI_DATA <= x"0" & CH5_1_rc;
            when 16#2F# => SPI_DATA <= x"0" & CH6_0_rc;
            when 16#30# => SPI_DATA <= x"0" & CH6_1_rc;
            when 16#31# => SPI_DATA <= x"0" & CH7_0_rc;
            when 16#32# => SPI_DATA <= x"0" & CH7_1_rc;
            when 16#33# => SPI_DATA <= x"0" & CH8_0_rc;
            when 16#34# => SPI_DATA <= x"0" & CH8_1_rc;
            when 16#35# => SPI_DATA <= x"0" & CH9_0_rc;
            when 16#36# => SPI_DATA <= x"0" & CH9_1_rc;
            when 16#37# => SPI_DATA <= x"0" & CH10_0_rc;
            when 16#38# => SPI_DATA <= x"0" & CH10_1_rc;
            when 16#39# => SPI_DATA <= x"0" & CH11_0_rc;
            when 16#3A# => SPI_DATA <= x"0" & CH11_1_rc;
            when 16#3B# => SPI_DATA <= x"0" & CH12_0_rc;
            when 16#3C# => SPI_DATA <= x"0" & CH12_1_rc;
            when 16#3D# => SPI_DATA <= x"0" & Ampl_sat;

            when 16#3E# => SPI_DATA <= pshift2(5) & pshift2(5) & pshift2 & pshift1(5) & pshift1(5) & pshift1;
            when 16#3F# => SPI_DATA <= x"00" & pshift3(5) & pshift3(5) & pshift3;

            when 16#40# => SPI_DATA <= "00" & TDC1A_raw (12 downto 7) & '0' & TDC1A_raw(6 downto 0);
            when 16#41# => SPI_DATA <= "00" & TDC1B_raw (12 downto 7) & '0' & TDC1B_raw(6 downto 0);
            when 16#42# => SPI_DATA <= "00" & TDC1C_raw (12 downto 7) & '0' & TDC1C_raw(6 downto 0);
            when 16#43# => SPI_DATA <= "00" & TDC1D_raw (12 downto 7) & '0' & TDC1D_raw(6 downto 0);
            when 16#44# => SPI_DATA <= "00" & TDC2A_raw (12 downto 7) & '0' & TDC2A_raw(6 downto 0);
            when 16#45# => SPI_DATA <= "00" & TDC2B_raw (12 downto 7) & '0' & TDC2B_raw(6 downto 0);
            when 16#46# => SPI_DATA <= "00" & TDC2C_raw (12 downto 7) & '0' & TDC2C_raw(6 downto 0);
            when 16#47# => SPI_DATA <= "00" & TDC2D_raw (12 downto 7) & '0' & TDC2D_raw(6 downto 0);
            when 16#48# => SPI_DATA <= "00" & TDC3A_raw (12 downto 7) & '0' & TDC3A_raw(6 downto 0);
            when 16#49# => SPI_DATA <= "00" & TDC3B_raw (12 downto 7) & '0' & TDC3B_raw(6 downto 0);
            when 16#4A# => SPI_DATA <= "00" & TDC3C_raw (12 downto 7) & '0' & TDC3C_raw(6 downto 0);
            when 16#4B# => SPI_DATA <= "00" & TDC3D_raw (12 downto 7) & '0' & TDC3D_raw(6 downto 0);

            when 16#4C# => SPI_DATA <= CH1_Z0;
            when 16#4D# => SPI_DATA <= CH1_Z1;
            when 16#4E# => SPI_DATA <= CH2_Z0;
            when 16#4F# => SPI_DATA <= CH2_Z1;
            when 16#50# => SPI_DATA <= CH3_Z0;
            when 16#51# => SPI_DATA <= CH3_Z1;
            when 16#52# => SPI_DATA <= CH4_Z0;
            when 16#53# => SPI_DATA <= CH4_Z1;
            when 16#54# => SPI_DATA <= CH5_Z0;
            when 16#55# => SPI_DATA <= CH5_Z1;
            when 16#56# => SPI_DATA <= CH6_Z0;
            when 16#57# => SPI_DATA <= CH6_Z1;
            when 16#58# => SPI_DATA <= CH7_Z0;
            when 16#59# => SPI_DATA <= CH7_Z1;
            when 16#5A# => SPI_DATA <= CH8_Z0;
            when 16#5B# => SPI_DATA <= CH8_Z1;
            when 16#5C# => SPI_DATA <= CH9_Z0;
            when 16#5D# => SPI_DATA <= CH9_Z1;
            when 16#5E# => SPI_DATA <= CH10_Z0;
            when 16#5F# => SPI_DATA <= CH10_Z1;
            when 16#60# => SPI_DATA <= CH11_Z0;
            when 16#61# => SPI_DATA <= CH11_Z1;
            when 16#62# => SPI_DATA <= CH12_Z0;
            when 16#63# => SPI_DATA <= CH12_Z1;

            when 16#64# => SPI_DATA <= std_logic_vector(resize(signed(CH1_0_rg), 16));
            when 16#65# => SPI_DATA <= std_logic_vector(resize(signed(CH1_1_rg), 16));
            when 16#66# => SPI_DATA <= std_logic_vector(resize(signed(CH2_0_rg), 16));
            when 16#67# => SPI_DATA <= std_logic_vector(resize(signed(CH2_1_rg), 16));
            when 16#68# => SPI_DATA <= std_logic_vector(resize(signed(CH3_0_rg), 16));
            when 16#69# => SPI_DATA <= std_logic_vector(resize(signed(CH3_1_rg), 16));
            when 16#6A# => SPI_DATA <= std_logic_vector(resize(signed(CH4_0_rg), 16));
            when 16#6B# => SPI_DATA <= std_logic_vector(resize(signed(CH4_1_rg), 16));
            when 16#6C# => SPI_DATA <= std_logic_vector(resize(signed(CH5_0_rg), 16));
            when 16#6D# => SPI_DATA <= std_logic_vector(resize(signed(CH5_1_rg), 16));
            when 16#6E# => SPI_DATA <= std_logic_vector(resize(signed(CH6_0_rg), 16));
            when 16#6F# => SPI_DATA <= std_logic_vector(resize(signed(CH6_1_rg), 16));
            when 16#70# => SPI_DATA <= std_logic_vector(resize(signed(CH7_0_rg), 16));
            when 16#71# => SPI_DATA <= std_logic_vector(resize(signed(CH7_1_rg), 16));
            when 16#72# => SPI_DATA <= std_logic_vector(resize(signed(CH8_0_rg), 16));
            when 16#73# => SPI_DATA <= std_logic_vector(resize(signed(CH8_1_rg), 16));
            when 16#74# => SPI_DATA <= std_logic_vector(resize(signed(CH9_0_rg), 16));
            when 16#75# => SPI_DATA <= std_logic_vector(resize(signed(CH9_1_rg), 16));
            when 16#76# => SPI_DATA <= std_logic_vector(resize(signed(CH10_0_rg), 16));
            when 16#77# => SPI_DATA <= std_logic_vector(resize(signed(CH10_1_rg), 16));
            when 16#78# => SPI_DATA <= std_logic_vector(resize(signed(CH11_0_rg), 16));
            when 16#79# => SPI_DATA <= std_logic_vector(resize(signed(CH11_1_rg), 16));
            when 16#7A# => SPI_DATA <= std_logic_vector(resize(signed(CH12_0_rg), 16));
            when 16#7B# => SPI_DATA <= std_logic_vector(resize(signed(CH12_1_rg), 16));

            when 16#7C# => SPI_DATA <= x"0" & chans_ena_r;
            when 16#7D# => SPI_DATA <= x"0" & Z_alarm;

            when 16#7F#           => SPI_DATA           <= x"0" & "00" & dcs_irq & BC_JUMP3 & BC_JUMP2 & BC_JUMP1 & GBTRXerr & GBTRX_ready & lock300_3 & lock300_2 & lock300_1 & lock320;
            when 16#80# to 16#BF# => SPI_DATA <= spi_buf_out;
            when 16#C0# to 16#EF# => SPI_DATA <= cnt_out;
            when 16#F0#           => SPI_DATA           <= rd_buf_vector(15 downto 0);
            when 16#F1#           => SPI_DATA           <= rd_buf_vector(31 downto 16);
            when 16#F2#           => SPI_DATA           <= rd_buf_vector(47 downto 32);
            when 16#F3#           => SPI_DATA           <= x"0" & rd_buf_vector(59 downto 48);

            when others => SPI_DATA <= x"0000";

          end case;
        else
          SPI_DATA <= SPI_DATA(14 downto 0) & MOSII;
        end if;

      end if;
    end if;
  end process;

  hspid_w32 <= hspi_wr_data & hspi_wr_data_l;

  wr_hspi32 <= '1' when (reg32_wr2 = '0') and (reg32_wr1 = '1') else
    '0';
  rd_hspi32 <= '1' when (reg32_rd2 = '0') and (reg32_rd1 = '1') else
    '0';
  str_reg32 <= '1' when (reg32_str2 = '0') and (reg32_str1 = '1') else
    '0';

  reg_wr_data <= spi_wr_data when (spi_wr_req = '1') else
    hspi_wr_data;
  reg_wr_addr <= spi_addr when (spi_wr_req = '1') else
    hspi_addr;

  err_report_fifo_rden <= '1' when (str_reg32 = '1') and (to_integer(unsigned(hspi_addr(7 downto 0))) = 16#F2#) else
    '0';
  readout_err_rden <= '1' when (str_reg32 = '1') and (to_integer(unsigned(hspi_addr(7 downto 0))) = 16#EA#) else
    '0';

  process (TX_CLK, sreset)
  begin
    if sreset = '1' then
      buf_vector   <= x"000000000000000";
      buf_cou      <= x"A0";
      dcs_irq      <= '0';
      vect_clr_req <= '0';
    else
      if (TX_CLK'event and TX_CLK = '1') then

        reg32_wr2   <= reg32_wr1;
        reg32_wr1   <= reg32_wr0;
        reg32_wr0   <= reg32_wr;
        reg32_rd2   <= reg32_rd1;
        reg32_rd1   <= reg32_rd0;
        reg32_rd0   <= reg32_rd;
        reg32_str2  <= reg32_str1;
        reg32_str1  <= reg32_str0;
        reg32_str0  <= reg32_str;
        spibuf_wr2  <= spibuf_wr1;
        spibuf_wr1  <= spibuf_wr0;
        spibuf_wr0  <= spibuf_wr;
        hspibuf_wr2 <= hspibuf_wr1;
        hspibuf_wr1 <= hspibuf_wr0;
        hspibuf_wr0 <= hspibuf_wr;
        spibuf_rd2  <= spibuf_rd1;
        spibuf_rd1  <= spibuf_rd0;
        spibuf_rd0  <= spibuf_rd;
        hspibuf_rd2 <= hspibuf_rd1;
        hspibuf_rd1 <= hspibuf_rd0;
        hspibuf_rd0 <= hspibuf_rd;

        buf_lock2 <= buf_lock1;
        buf_lock1 <= buf_lock0;
        buf_lock0 <= buf_lock;

        hbuf_req <= (not hspibuf_wr2) and hspibuf_wr1 and sbuf_wrena;

        --err_report_fifo_rden <= '0';
        if (rd_hspi32 = '1') then

          if (rdo_sel = '1') then
            hspib_32 <= ipbus_status_reg(to_integer(unsigned(hspi_addr(7 downto 0))) - 16#E8#);
            --if (to_integer(unsigned(hspi_addr(7 downto 0)))-16#E8#) = 10 then err_report_fifo_rden <= '1';  end if;
          else
            if (flsh_sel = '1') then
              hspib_32 <= hspid_r32;
            end if;

          end if;
        end if;
        if (hbuf_wrena = '1') and (hspi_addr(5 downto 0) < "111100") then
          buf_vector(to_integer(unsigned(hspi_addr(5 downto 0)))) <= '1';
          buf_cou                                                 <= x"00";
          if (vect_clr = '1') then
            vect_clr_req <= '1';
          end if;
        else
          vect_clr_req <= '0';
          if (vect_clr = '1') or (vect_clr_req = '1') then
            rd_buf_vector <= buf_vector;
            buf_vector    <= x"000000000000000";
          end if;
          if (buf_cou /= x"A0") then
            buf_cou <= buf_cou + 1;
          end if;

        end if;
        if (buf_cou = x"9F") then
          dcs_irq <= '1';
        else
          if (stat_clr1 = '1') and (stat_clr = '0') then
            dcs_irq <= '0';
          end if;
        end if;

        if (reg32_wr2 = '0') and (reg32_wr1 = '1') and (hspi_addr(7 downto 0) <= 16#E7#) then
          if (hspi_addr(7 downto 0) = 16#D8#) then
            ipbus_control_reg(0) <= hspid_w32;
          else
            ipbus_control_reg(to_integer(unsigned(hspi_addr(7 downto 0))) - 16#D8#) <= hspid_w32;
          end if;
        end if;

      end if;
    end if;
  end process;

  vect_clr   <= (not buf_lock2) and buf_lock1;
  sbuf_wrena <= (not spibuf_wr2) and spibuf_wr1;
  sbuf_rdena <= (not spibuf_rd2) and spibuf_rd1;
  hbuf_wrena <= ((not hspibuf_wr2) and hspibuf_wr1 and (not sbuf_wrena)) or hbuf_req;
  hbuf_rdena <= (not hspibuf_rd2) and hspibuf_rd1;
  sbuf_ena   <= sbuf_wrena or sbuf_rdena;
  hbuf_ena   <= hbuf_wrena or hbuf_rdena;

  Xmegamem : Xmega_buf port
  map (clka => TX_CLK, ena => hbuf_ena, wea(0) => hbuf_wrena, addra => hspi_addr(5 downto 0), dina => hspi_wr_data, douta => hspi_buf_out, clkb => TX_CLK, enb => sbuf_ena, web(0) => sbuf_wrena, addrb => spi_addr(5 downto 0), dinb => spi_wr_data, doutb => spi_buf_out);

  tcm_req <= ((not tcm_req2) and tcm_req1) or ((not gs0_1) and gs0_0) or ((not gs1_1) and gs1_0);

  reg32_320_wr  <= reg32_320_wr1 and (not reg32_320_wr2);
  reg32_320_str <= reg32_320_str1 and (not reg32_320_str2);

  process (clk320)
  begin
    if (clk320'event and clk320 = '1') then

      reg32_320_wr2  <= reg32_320_wr1;
      reg32_320_wr1  <= reg32_320_wr0;
      reg32_320_wr0  <= reg32_wr;
      reg32_320_str2 <= reg32_320_str1;
      reg32_320_str1 <= reg32_320_str0;
      reg32_320_str0 <= reg32_str;

      gs0_1 <= gs0_0;
      gs0_0 <= gbt_global_status(0);
      gs1_1 <= gs1_0;
      gs1_0 <= gbt_global_status(1);

      spi_wr2  <= spi_wr1;
      spi_wr1  <= spi_wr0;
      spi_wr0  <= spi_wr_rdy;
      hspi_wr2 <= hspi_wr1;
      hspi_wr1 <= hspi_wr0;
      hspi_wr0 <= hspi_wr_rdy;

      tcm_req2 <= tcm_req1;
      tcm_req1 <= tcm_req0;
      tcm_req0 <= tcm_reqh;

      if (spi_wr2 = '0') and (spi_wr1 = '1') then
        spi_wr_req <= '1';
      end if;
      if (hspi_wr2 = '0') and (hspi_wr1 = '1') then
        hspi_wr_req <= '1';
      end if;

      if (cnt_rst = '1') then
        cnt_rst <= '0';
      end if;
      if (hyst_rst = '1') then
        hyst_rst <= '0';
      end if;

      if (sreset = '1') then
        chans_block <= '0';
        hyst_md(15) <= '0';
        is_rst      <= '1';
      else
        if (spi_wr_req = '1') or (hspi_wr_req = '1') then
          case reg_wr_addr(7 downto 0) is
            when x"00" => gate_time_high <= reg_wr_data(7 downto 0);
              if (spi_wr_req = '0') then
                fdd <= reg_wr_data(8);
              end if;
            when x"01" => CH1A_shift <= reg_wr_data(11 downto 0);
              if (spi_wr_req = '0') then
                trig_dis(0) <= reg_wr_data(12);
              end if;
            when x"02" => CH1B_shift <= reg_wr_data(11 downto 0);
              if (spi_wr_req = '0') then
                trig_dis(1) <= reg_wr_data(12);
              end if;
            when x"03" => CH1C_shift <= reg_wr_data(11 downto 0);
              if (spi_wr_req = '0') then
                trig_dis(2) <= reg_wr_data(12);
              end if;
            when x"04" => CH1D_shift <= reg_wr_data(11 downto 0);
              if (spi_wr_req = '0') then
                trig_dis(3) <= reg_wr_data(12);
              end if;
            when x"05" => CH2A_shift <= reg_wr_data(11 downto 0);
              if (spi_wr_req = '0') then
                trig_dis(4) <= reg_wr_data(12);
              end if;
            when x"06" => CH2B_shift <= reg_wr_data(11 downto 0);
              if (spi_wr_req = '0') then
                trig_dis(5) <= reg_wr_data(12);
              end if;
            when x"07" => CH2C_shift <= reg_wr_data(11 downto 0);
              if (spi_wr_req = '0') then
                trig_dis(6) <= reg_wr_data(12);
              end if;
            when x"08" => CH2D_shift <= reg_wr_data(11 downto 0);
              if (spi_wr_req = '0') then
                trig_dis(7) <= reg_wr_data(12);
              end if;
            when x"09" => CH3A_shift <= reg_wr_data(11 downto 0);
              if (spi_wr_req = '0') then
                trig_dis(8) <= reg_wr_data(12);
              end if;
            when x"0A" => CH3B_shift <= reg_wr_data(11 downto 0);
              if (spi_wr_req = '0') then
                trig_dis(9) <= reg_wr_data(12);
              end if;
            when x"0B" => CH3C_shift <= reg_wr_data(11 downto 0);
              if (spi_wr_req = '0') then
                trig_dis(10) <= reg_wr_data(12);
              end if;
            when x"0C" => CH3D_shift <= reg_wr_data(11 downto 0);
              if (spi_wr_req = '0') then
                trig_dis(11) <= reg_wr_data(12);
              end if;
            when x"25" => CH1_0_rc  <= reg_wr_data(11 downto 0);
            when x"26" => CH1_1_rc  <= reg_wr_data(11 downto 0);
            when x"27" => CH2_0_rc  <= reg_wr_data(11 downto 0);
            when x"28" => CH2_1_rc  <= reg_wr_data(11 downto 0);
            when x"29" => CH3_0_rc  <= reg_wr_data(11 downto 0);
            when x"2A" => CH3_1_rc  <= reg_wr_data(11 downto 0);
            when x"2B" => CH4_0_rc  <= reg_wr_data(11 downto 0);
            when x"2C" => CH4_1_rc  <= reg_wr_data(11 downto 0);
            when x"2D" => CH5_0_rc  <= reg_wr_data(11 downto 0);
            when x"2E" => CH5_1_rc  <= reg_wr_data(11 downto 0);
            when x"2F" => CH6_0_rc  <= reg_wr_data(11 downto 0);
            when x"30" => CH6_1_rc  <= reg_wr_data(11 downto 0);
            when x"31" => CH7_0_rc  <= reg_wr_data(11 downto 0);
            when x"32" => CH7_1_rc  <= reg_wr_data(11 downto 0);
            when x"33" => CH8_0_rc  <= reg_wr_data(11 downto 0);
            when x"34" => CH8_1_rc  <= reg_wr_data(11 downto 0);
            when x"35" => CH9_0_rc  <= reg_wr_data(11 downto 0);
            when x"36" => CH9_1_rc  <= reg_wr_data(11 downto 0);
            when x"37" => CH10_0_rc <= reg_wr_data(11 downto 0);
            when x"38" => CH10_1_rc <= reg_wr_data(11 downto 0);
            when x"39" => CH11_0_rc <= reg_wr_data(11 downto 0);
            when x"3A" => CH11_1_rc <= reg_wr_data(11 downto 0);
            when x"3B" => CH12_0_rc <= reg_wr_data(11 downto 0);
            when x"3C" => CH12_1_rc <= reg_wr_data(11 downto 0);
            when x"3D" => Ampl_sat  <= reg_wr_data(11 downto 0);
              ampl_low                <= reg_wr_data(15 downto 12);

            when x"7C" => chans_ena_r <= reg_wr_data(11 downto 0);

            when x"7E" => hyst_md(14 downto 0) <= reg_wr_data(14) & '0' & reg_wr_data(12 downto 0);
              if (hyst_rst = '0') and (reg_wr_data(13) = '1') then
                hyst_rst <= '1';
              end if;

            when x"7F" =>
              if (cnt_rst = '0') and (reg_wr_data(9) = '1') then
                cnt_rst <= '1';
              end if;
              if (hspi_wr_req = '1') and (spi_wr_req = '0') then
                cnt_md <= reg_wr_data(10);
              end if;
              if (hspi_wr_req = '1') and (spi_wr_req = '0') and (reg_wr_data(11) = '1') then
                is_rst <= '0';
              end if;
              if (spi_wr_req = '1') and (reg_wr_data(11) = '1') then
                chans_block <= '1';
              end if;

            when others => null;
          end case;
          if (spi_wr_req = '1') then
            spi_wr_req <= '0';
          end if;
          if (hspi_wr_req = '1') and (spi_wr_req = '0') then
            hspi_wr_req <= '0';
          end if;

        end if;
        if ((spi_wr_req = '1') or (hspi_wr_req = '1')) and (reg_wr_addr(7 downto 0) = x"7E") then
          hyst_md(15) <= reg_wr_data(15);
        else
          if (hyst_stp = '1') then
            hyst_md(15) <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;

  RESET     <= not rsti;
  spi_rden  <= SPI_CS;
  hspi_rden <= not HSELI;

  HMISOI <= HSPI_DATA(15);

  gate_time_low <= (not gate_time_high) + 1;

  rd_lock <= rd_lock_spi or rd_lock_hspi;

  ch_en : for i in 0 to 11 generate

    chans_ena(i) <= chans_ena_r(i) and chans_block;

  end generate;

  process (tdcclk1)
  begin
    if (tdcclk1'event and tdcclk1 = '1') then

      spi_lock_1  <= spi_lock0_1;
      spi_lock0_1 <= rd_lock;

    end if;
  end process;

  process (tdcclk2)
  begin
    if (tdcclk2'event and tdcclk2 = '1') then

      spi_lock_2  <= spi_lock0_2;
      spi_lock0_2 <= rd_lock;

    end if;
  end process;

  process (tdcclk3)
  begin
    if (tdcclk3'event and tdcclk3 = '1') then

      spi_lock_3  <= spi_lock0_3;
      spi_lock0_3 <= rd_lock;

    end if;
  end process;

  process (clk300_1)
  begin
    if (clk300_1'event and clk300_1 = '1') then

      almclr10 <= ALM_CLR;
      almclr11 <= almclr10;
      alm_clr1 <= almclr11;
      hclr10   <= Hs_rd;
      hclr11   <= hclr10;
      h_clr1   <= hclr11;

      BC_STR11 <= BC_STR1;
      BC_STR12 <= BC_STR11;

      TDC_COU1 <= TDC_COU1 + 1;

      if (BC_STR1 = '1' and BC_STR11 = '0') then
        BC_PER1 <= TDC_COU1 & BC_BITS1;
      end if;

      if (BC_STR11 = '1' and BC_STR12 = '0') then
        BCOLD1 <= BC_PER1(1 downto 0);
      end if;

      if (BC_STR11 = '1' and BC_STR12 = '0') and (BCOLD1 /= BC_PER1(1 downto 0)) then
        BC_JUMP1  <= '1';
        HBC_JUMP1 <= '1';
        jumpa1    <= '1';
      else
        jumpa1 <= '0';
        if (alm_clr1 = '0') and (almclr11 = '1') then
          BC_JUMP1 <= '0';
        end if;
        if (h_clr1 = '0') and (hclr11 = '1') then
          HBC_JUMP1 <= '0';
        end if;
      end if;

    end if;
  end process;

  process (clk300_2)
  begin
    if (clk300_2'event and clk300_2 = '1') then

      almclr20 <= ALM_CLR;
      almclr21 <= almclr20;
      alm_clr2 <= almclr21;
      hclr20   <= Hs_rd;
      hclr21   <= hclr20;
      h_clr2   <= hclr21;

      BC_STR21 <= BC_STR2;
      BC_STR22 <= BC_STR21;

      TDC_COU2 <= TDC_COU2 + 1;

      if (BC_STR2 = '1' and BC_STR21 = '0') then
        BC_PER2 <= TDC_COU2 & BC_BITS2;
      end if;
      if (BC_STR21 = '1' and BC_STR22 = '0') then
        BCOLD2 <= BC_PER2(1 downto 0);
      end if;
      if BC_STR21 = '1' and BC_STR22 = '0' and (BCOLD2 /= BC_PER2(1 downto 0)) then
        BC_JUMP2  <= '1';
        HBC_JUMP2 <= '1';
        jumpa2    <= '1';
      else
        jumpa2 <= '0';
        if (alm_clr2 = '0') and (almclr21 = '1') then
          BC_JUMP2 <= '0';
        end if;
        if (h_clr2 = '0') and (hclr21 = '1') then
          HBC_JUMP2 <= '0';
        end if;
      end if;

    end if;
  end process;

  process (clk300_3)
  begin
    if (clk300_3'event and clk300_3 = '1') then

      almclr30 <= ALM_CLR;
      almclr31 <= almclr30;
      alm_clr3 <= almclr31;
      hclr30   <= Hs_rd;
      hclr31   <= hclr30;
      h_clr3   <= hclr31;

      BC_STR31 <= BC_STR3;
      BC_STR32 <= BC_STR31;

      TDC_COU3 <= TDC_COU3 + 1;

      if (BC_STR3 = '1' and BC_STR31 = '0') then
        BC_PER3 <= TDC_COU3 & BC_BITS3;
      end if;
      if (BC_STR31 = '1' and BC_STR32 = '0') then
        BCOLD3 <= BC_PER3(1 downto 0);
      end if;
      if BC_STR31 = '1' and BC_STR32 = '0' and (BCOLD3 /= BC_PER3(1 downto 0)) then
        BC_JUMP3  <= '1';
        HBC_JUMP3 <= '1';
        jumpa3    <= '1';
      else
        jumpa3 <= '0';
        if (alm_clr3 = '0') and (almclr31 = '1') then
          BC_JUMP3 <= '0';
        end if;
        if (h_clr3 = '0') and (hclr31 = '1') then
          HBC_JUMP3 <= '0';
        end if;
      end if;

    end if;
  end process;

  PM_data_toreadout.data_word <= data_word;
  process (clk320)
  begin
    if (clk320'event and clk320 = '1') then

      rx_phase_status(2 downto 0) <= readout_status.rx_phase;
      rx_phase_status(3)          <= readout_status.Rx_Phase_error;

      spi_lock320    <= spi_lock320_0;
      spi_lock320_0  <= rd_lock;
      hspi_lock320   <= hspi_lock320_0;
      hspi_lock320_0 <= rd_lock_hspi;
      tto            <= tt;
      tao            <= ta;
      MCLK40_0       <= MCLK40T;
      MCLK40_1       <= MCLK40_0;
      if (MCLK40_0 /= MCLK40_1) then
        mt_cou <= "000";
      else
        mt_cou <= mt_cou + 1;
      end if;

      PM_data_toreadout.is_header <= is_header;
      is_header                   <= wr_out_id;
      PM_data_toreadout.is_data   <= is_data;
      is_data                     <= Event_ready or wr_out_id;
      data_word                   <= DATA80_in;

      if (wr_out_id = '1') then
        DATA80_in <= x"F" & '0' & WRDS_NUM & x"000000" & rx_phase_status & EV_ID_out(55 downto 12);
      else
        DATA80_in <= EV_DATA80;
      end if;
      if (Event_free = '1') or (wr_out_id = '1') then
        ev_tout_cnt <= (others => '0');
      else
        ev_tout_cnt <= ev_tout_cnt + 1;
      end if;
      if (ev_tout_cnt = 96) and (wr_out_id = '0') then
        ev_tout <= '1';
      else
        ev_tout <= '0';
      end if;
      ev_tout0 <= ev_tout;

      --if (wr_out_id='1') or (Event_ready='1') then WR_fifo_out<='1'; else WR_fifo_out<='0';  end if;

      if (Event_ready = '0') then
        if (Event_ready_0 = '1') and (ev_tout = '0') then
          Event_ready <= '1';
        end if;
      else
        if (CH_do = 0) then
          Event_ready <= '0';
        end if;
      end if;
      if (wr_nch = '1') then
        CH_do  <= EV_ID_out(11 downto 0);
        wr_nch <= '0';
      else
        if (Event_ready = '1') or (Event_ready_0 = '1') then

          case CH_N0_0 is
            when x"1"   => CH_do(0)  <= '0';
            when x"2"   => CH_do(1)  <= '0';
            when x"3"   => CH_do(2)  <= '0';
            when x"4"   => CH_do(3)  <= '0';
            when x"5"   => CH_do(4)  <= '0';
            when x"6"   => CH_do(5)  <= '0';
            when x"7"   => CH_do(6)  <= '0';
            when x"8"   => CH_do(7)  <= '0';
            when x"9"   => CH_do(8)  <= '0';
            when x"A"   => CH_do(9)  <= '0';
            when x"B"   => CH_do(10) <= '0';
            when x"C"   => CH_do(11) <= '0';
            when others => null;
          end case;

          case CH_N1_0 is
            when x"2"   => CH_do(1)  <= '0';
            when x"3"   => CH_do(2)  <= '0';
            when x"4"   => CH_do(3)  <= '0';
            when x"5"   => CH_do(4)  <= '0';
            when x"6"   => CH_do(5)  <= '0';
            when x"7"   => CH_do(6)  <= '0';
            when x"8"   => CH_do(7)  <= '0';
            when x"9"   => CH_do(8)  <= '0';
            when x"A"   => CH_do(9)  <= '0';
            when x"B"   => CH_do(10) <= '0';
            when x"C"   => CH_do(11) <= '0';
            when others => null;
          end case;
        end if;
        if (sreset = '0') and (EV_ID_rd = '1') then
          wr_nch <= '1';
        end if;
      end if;

      if (sreset = '1') then
        Event_free <= '1';
      else
        if (Event_free = '1') then
          if (EV_ID_empty = '0') then
            EVENT_free <= '0';
          end if;
        else
          if (((Event_ready = '1') and (CH_do = 0)) or (ev_tout0 = '1')) and (EV_ID_empty = '1') then
            Event_free <= '1';
          end if;
        end if;
      end if;

      if (Event_ready = '1') or (Event_ready_0 = '1') then
        CH_N0 <= CH_N0_0;
        CH_N1 <= CH_N1_0;
      end if;

      if (mt_cou = "001") then
        if (New_BCID = '1') then
          BC_COU   <= readout_status. BCID_from_CRU_corrected;
          Orbit_ID <= readout_status. ORBIT_from_CRU_corrected;
          if (readout_status. BCID_from_CRU_corrected > x"003") then
            TR_to <= readout_status. BCID_from_CRU_corrected(5 downto 0) - "000100";
          else
            TR_to <= "1010" & readout_status. BCID_from_CRU_corrected(1 downto 0);
          end if;

        else
          if (BC_COU = x"DEB") then
            BC_cou   <= x"000";
            Orbit_ID <= Orbit_ID + 1;
          else
            BC_cou <= BC_cou + 1;
          end if;
          if (BC_COU > x"003") then
            TR_to <= BC_COU(5 downto 0) - "000100";
          else
            TR_to <= "1010" & BC_COU(1 downto 0);
          end if;
        end if;
      end if;

      if ((EV_ID_out(23 downto 12) = hyst_md(11 downto 0)) or (hyst_md(12) = '0')) and (hyst_md(15) = '1') then
        start_hyst <= Event_ready_0 and (not Event_ready);
      else
        start_hyst <= '0';
      end if;
    end if;
  end process;

  New_BCID <= readout_status.bc_delay_apply;

  CH_N0_0 <= x"1" when CH_do(0) = '1'
    else
    x"2" when CH_do(1) = '1'
    else
    x"3" when CH_do(2) = '1'
    else
    x"4" when CH_do(3) = '1'
    else
    x"5" when CH_do(4) = '1'
    else
    x"6" when CH_do(5) = '1'
    else
    x"7" when CH_do(6) = '1'
    else
    x"8" when CH_do(7) = '1'
    else
    x"9" when CH_do(8) = '1'
    else
    x"A" when CH_do(9) = '1'
    else
    x"B" when CH_do(10) = '1'
    else
    x"C" when CH_do(11) = '1'
    else
    x"0";

  CH_N1_0 <= x"2" when CH_do(1) = '1' and (CH_N0_0 /= x"2")
    else
    x"3" when CH_do(2) = '1' and (CH_N0_0 /= x"3")
    else
    x"4" when CH_do(3) = '1' and (CH_N0_0 /= x"4")
    else
    x"5" when CH_do(4) = '1' and (CH_N0_0 /= x"5")
    else
    x"6" when CH_do(5) = '1' and (CH_N0_0 /= x"6")
    else
    x"7" when CH_do(6) = '1' and (CH_N0_0 /= x"7")
    else
    x"8" when CH_do(7) = '1' and (CH_N0_0 /= x"8")
    else
    x"9" when CH_do(8) = '1' and (CH_N0_0 /= x"9")
    else
    x"A" when CH_do(9) = '1' and (CH_N0_0 /= x"A")
    else
    x"B" when CH_do(10) = '1' and (CH_N0_0 /= x"B")
    else
    x"C" when CH_do(11) = '1' and (CH_N0_0 /= x"C")
    else
    x"0";
  EV_DATA80(32 downto 0) <= Data_out(0) when CH_N0 = x"1" else
  Data_out(1) when CH_N0 = x"2" else
  Data_out(2) when CH_N0 = x"3" else
  Data_out(3) when CH_N0 = x"4" else
  Data_out(4) when CH_N0 = x"5" else
  Data_out(5) when CH_N0 = x"6" else
  Data_out(6) when CH_N0 = x"7" else
  Data_out(7) when CH_N0 = x"8" else
  Data_out(8) when CH_N0 = x"9" else
  Data_out(9) when CH_N0 = x"A" else
  Data_out(10) when CH_N0 = x"B" else
  Data_out(11) when CH_N0 = x"C" else
  "0" & x"00000000";

  EV_DATA80(35 downto 33) <= "000";
  EV_DATA80(39 downto 36) <= CH_N0;

  EV_DATA80(72 downto 40) <= Data_out(1) when CH_N1 = x"2" else
  Data_out(2) when CH_N1 = x"3" else
  Data_out(3) when CH_N1 = x"4" else
  Data_out(4) when CH_N1 = x"5" else
  Data_out(5) when CH_N1 = x"6" else
  Data_out(6) when CH_N1 = x"7" else
  Data_out(7) when CH_N1 = x"8" else
  Data_out(8) when CH_N1 = x"9" else
  Data_out(9) when CH_N1 = x"A" else
  Data_out(10) when CH_N1 = x"B" else
  Data_out(11) when CH_N1 = x"C" else
  "0" & x"00000000";

  EV_DATA80(75 downto 73) <= "000";
  EV_DATA80(79 downto 76) <= CH_N1;
  inp_event               <= Event_in(0) or Event_in(1) or Event_in(2) or Event_in(3) or Event_in(4) or Event_in(5) or Event_in(6) or Event_in(7) or Event_in(8) or Event_in(9) or Event_in(10) or Event_in(11);
  Event_ready_0           <= ((not EV_ID_out(0)) or Data_rdy(0)) and ((not EV_ID_out(1)) or Data_rdy(1)) and ((not EV_ID_out(2)) or Data_rdy(2)) and ((not EV_ID_out(3)) or Data_rdy(3)) and ((not EV_ID_out(4)) or Data_rdy(4)) and ((not EV_ID_out(5)) or Data_rdy(5))
    and ((not EV_ID_out(6)) or Data_rdy(6)) and ((not EV_ID_out(7)) or Data_rdy(7)) and ((not EV_ID_out(8)) or Data_rdy(8)) and ((not EV_ID_out(9)) or Data_rdy(9)) and ((not EV_ID_out(10)) or Data_rdy(10)) and ((not EV_ID_out(11)) or Data_rdy(11))
    and not (Event_free or wr_nch);
  CH_NUM1  <= ("00" & EV_ID_out(0)) + ("00" & EV_ID_out(1)) + ("00" & EV_ID_out(2)) + ("00" & EV_ID_out(3)) + ("00" & EV_ID_out(4)) + ("00" & EV_ID_out(5));
  CH_NUM2  <= ("00" & EV_ID_out(6)) + ("00" & EV_ID_out(7)) + ("00" & EV_ID_out(8)) + ("00" & EV_ID_out(9)) + ("00" & EV_ID_out(10)) + ("00" & EV_ID_out(11));
  CH_NUM   <= ('0' & CH_NUM1) + ('0' & CH_NUM2);
  WRDS_NUM <= CH_NUM(3 downto 1) + ("00" & CH_NUM(0)) when (ev_tout = '0') else
    "000";

  FIFO_RD : for i in 0 to 11 generate
    DATA_rd(i) <= '1' when (Event_Ready_0 = '1') and (Event_Ready = '0') and (EV_ID_out(i) = '1') and (Data_rdy(i) = '1') else
    '0';
  end generate;

  FIFO_dis  <= EV_ID_empty and EVENT_free;
  wr_out_id <= (Event_ready_0 and (not Event_ready)) or ev_tout;

  --la2i(0)<=EVNTI; la2i(1)<=Zcal_done; la2i(2)<=inp_cou(1); la2i(3)<=CSTR2; la2i(4)<=inp_cou(2); la2i(5)<=CSTR3; la2i(6)<=inp_cou(3); la2i(7)<=CSTR4; la2i(8)<=inp_cou(4); la2i(9)<=CSTR5; la2i(10)<=inp_cou(5); la2i(11)<=CSTR6; 
  --la2i(12)<=inp_cou(6); la2i(13)<=CSTR7; la2i(14)<=inp_cou(7); la2i(15)<=CSTR8; lack2i<=inp_cou(8); lack3i<=CSTR9; la3i(14)<=inp_cou(9); la3i(15)<=CSTR10; la3i(12)<=inp_cou(10); la3i(13)<=CSTR11; la3i(10)<=inp_cou(11); la3i(11)<=CSTR12;

  --la2i(1 downto 0)<=BCOLD1(1 downto 0); la2i(2)<=BC_JUMP1; la2i(3)<=ALM_CLR; la2i(4)<=BC_JUMP2; la2i(5)<=BC_JUMP3;

  --la3i(0)<=rchange1; la3i(1)<=rchange2; la3i(2)<=rchange3;
  --la0i(0)<=MCLK40_IN1; la0i(1)<=MCLK40_IN2; la0i(2)<=MCLK40_IN3; la0i(3)<=CSTR1; la0i(4)<=CGE1; la0i(5)<=lTDCCLK1; la0i(6)<=RSA1;
  --la3i(15)<=inp_event;
  --la1i(15 downto 14) <= ttla;
  --la2i(15 downto 14) <= tala;

  --la2i(0)<=HSELI; la2i(1)<=HSCKI; la2i(2)<=HMOSII; la2i(3)<=HMISOI; la2i(4)<=hspi_h; la2i(5)<=rd_hyst_d0; la2i(6)<=hbuf_ena; la2i(7)<=hbuf_wrena; la2i(8)<=reg32_wr;

  --la3i(0)<=gs0;  la3i(1)<=gs1;
  --la2i(15) <= PM_data_toreadout.is_data;
  --la2i(14) <= PM_data_toreadout.is_packet;
  --la2i(13) <= PM_data_toreadout.is_header;
  --la2i(12 downto 0) <= PM_data_toreadout.data_word(12 downto 0);

end RTL;